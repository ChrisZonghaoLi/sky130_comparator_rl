** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp_tb.sch
**.subckt double_tail_comp_tb Di_n Di_p Vout_n Vout_p Q Q_bar Di_n_mc Di_p_mc Vout_n_mc Vout_p_mc
*+ Di_n_ms Di_p_ms Vout_n_ms Vout_p_ms Di_n_kn Di_p_kn Vout_n_kn Vout_p_kn
*.opin Di_n
*.opin Di_p
*.opin Vout_n
*.opin Vout_p
*.opin Q
*.opin Q_bar
*.opin Di_n_mc
*.opin Di_p_mc
*.opin Vout_n_mc
*.opin Vout_p_mc
*.opin Di_n_ms
*.opin Di_p_ms
*.opin Vout_n_ms
*.opin Vout_p_ms
*.opin Di_n_kn
*.opin Di_p_kn
*.opin Vout_n_kn
*.opin Vout_p_kn
x1 net1 Vclk_bar Vout_n Vout_p Di_n Di_p Vcm net10 Vclk GND double_tail_comp
VDD net1 net9 VDD
Vclk Vclk GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar Vclk_bar GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm Vcm GND dc Vcm
Vdiff net10 Vcm dc Vin
C2 Q_bar GND 10f m=1
C3 Q GND 10f m=1
x2 net17 Vout_n Q Vout_p Q_bar RS_latch
x3 net4 net3 Vout_n_mc Vout_p_mc Di_n_mc Di_p_mc net2 Vsc net15 GND double_tail_comp
VDD2 net4 GND VDD
Vclk2 net15 GND PULSE(0 VDD 0 Tr Tf Tclk_pk Tclk 0)
Vclk_bar2 net3 GND PULSE(0 VDD Tclk_pk Tr Tf Tclk_pk Tclk 0)
Vcm2 net2 GND dc Vcm
ASRC1 %v([ Vsc ]) filesrc
x4 net8 net7 Vout_n_ms Vout_p_ms Di_n_ms Di_p_ms net5 net6 net16 GND double_tail_comp
VDD3 net8 GND VDD
Vclk3 net16 GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar3 net7 GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm3 net5 GND dc Vcm
Vdiff2 net6 net5 dc Vin_min
VDD_latch net17 GND VDD
Rdummy net9 GND 1 m=1
x5 net13 net12 Vout_n_kn Vout_p_kn Di_n_kn Di_p_kn Vn_kn Vp_kn net18 GND double_tail_comp
VDD4 net13 GND VDD
Vclk4 net18 GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar5 net12 GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm4 net11 GND dc Vcm
Vdiff4 net14 net11 dc Vin
Rdummyn net11 Vn_kn 8k m=1
Rdummyp net14 Vp_kn 8k m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



*.OPTIONS maxord=1
*.OPTIONS itl1=200
*.OPTIONS itl2=200
*.OPTIONS itl4=200

* save all voltage and current
.save all
.options savecurrents
.options seed=random

.nodeset V(Vout_n) = 0
.nodeset V(Vout_p) = 0
.nodeset V(Di_n) = 0
.nodeset V(Di_p) = 0
.nodeset V(Q) = 0
.nodeset V(Q_bar) = 0

.nodeset V(Vout_n_mc) = 0
.nodeset V(Vout_p_mc) = 0
.nodeset V(Di_n_mc) = 0
.nodeset V(Di_p_mc) = 0

.nodeset V(Vout_n_ms) = 0
.nodeset V(Vout_p_ms) = 0
.nodeset V(Di_n_ms) = 0
.nodeset V(Di_p_ms) = 0

.control
set filetype=ascii
set units=degrees

.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/sky130_comparator/xschem/simulations/double_tail_comp_tb_vars.spice
.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/sky130_comparator/xschem/simulations/double_tail_comp_tb_analyses.spice

.endc


**** end user architecture code
**.ends

* expanding   symbol:  double_tail_comp.sym # of pins=10
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp.sch
.subckt double_tail_comp VDD CLK_bar Vout_n Vout_p Di_p Di_n Vin_n Vin_p CLK VSS
*.ipin CLK
*.ipin Vin_p
*.ipin Vin_n
*.opin Di_n
*.opin Di_p
*.opin Vout_n
*.opin Vout_p
*.ipin CLK_bar
*.iopin VDD
*.iopin VSS
XM1 Di_n Vin_p net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=W_M1 nf=10 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Di_p Vin_n net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=W_M2 nf=10 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Di_n CLK VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=W_M3 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Di_p CLK VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=W_M4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 CLK VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=W_M5 nf=12 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vout_p Di_n VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=W_M6 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout_p Vout_n VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=W_M7 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 Vout_n Vout_p VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=W_M8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 Vout_n Di_p VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=W_M9 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 Vout_p Vout_n net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=W_M10 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 Vout_n Vout_p net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=W_M11 nf=2 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net2 CLK_bar VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=W_M12 nf=12 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  RS_latch.sym # of pins=5
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/RS_latch.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/RS_latch.sch
.subckt RS_latch VDD R Q S Q_bar
*.iopin VDD
*.opin Q
*.opin Q_bar
*.ipin R
*.ipin S
x1 VDD R Q_bar Q nor
x2 VDD Q S Q_bar nor
.ends


* expanding   symbol:  nor.sym # of pins=4
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/nor.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/nor.sch
.subckt nor VDD A B out
*.iopin VDD
*.ipin A
*.ipin B
*.opin out
XM1 out B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out B net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
**** begin user architecture code

.model filesrc filesource (file="staircase_voltage.txt" amploffset=[Vcm] amplscale=[1] timeoffset=0
+ timescale=1 timerelative=false amplstep=false)

**** end user architecture code
.end

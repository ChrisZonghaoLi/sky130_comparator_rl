.param W_M1=5.5357814729213715
.param W_M3=4.901380236297846
.param W_M5=5.485002116709947
.param W_M6=9.855662246569992
.param W_M7=4.927831123284996
.param W_M10=5.436397657878697
.param W_M12=4.9983246502652765
.param W_M2=W_M1
.param W_M4=W_M3
.param W_M9=W_M6
.param W_M8=W_M7
.param W_M11=W_M10
.param Vcm=1.0474329798482358
.param VDD=1.8
.param Vin=0.05
.param Vin_min=0.0001
.param CL=2e-14
.param Tclk=1e-09
.param Tclk_pk=4.5e-10
.param Tdelay=2e-10
.param Tdelay_bar=7.000000000000001e-10
.param Tr=5.000000000000001e-11
.param Tf=5.000000000000001e-11

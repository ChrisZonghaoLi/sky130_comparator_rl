magic
tech sky130A
timestamp 1706848095
<< pwell >>
rect 0 0 144 504
<< end >>

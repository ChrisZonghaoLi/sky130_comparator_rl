.param W_M1=9.054640832543374e-06
.param W_M3=1.4282417398691177e-06
.param W_M5=3.6263448050618174e-06
.param W_M6=4.6464409351348867e-07
.param W_M7=2.3232204675674433e-07
.param W_M10=6.184994107484818e-07
.param W_M12=9.782913843393328e-06
.param W_M2=W_M1
.param W_M4=W_M3
.param W_M9=W_M6
.param W_M8=W_M7
.param W_M11=W_M10
.param Vcm=1.0666197180747985
.param VDD=3.3
.param Vin=0.05
.param Vin_min=0.0001
.param CL=2e-14
.param Tclk=1e-09
.param Tclk_pk=4.5e-10
.param Tdelay=2e-10
.param Tdelay_bar=7.000000000000001e-10
.param Tr=5.000000000000001e-11
.param Tf=5.000000000000001e-11

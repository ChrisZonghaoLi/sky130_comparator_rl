magic
tech sky130A
timestamp 1706848148
<< nwell >>
rect 0 0 144 504
<< end >>

magic
tech sky130A
timestamp 1704925934
<< checkpaint >>
rect -650 -660 3962 1668
<< metal1 >>
rect 1497 844 1527 1028
rect 1641 844 1671 1028
rect 1497 -20 1527 164
rect 1641 -20 1671 164
<< metal2 >>
rect -20 978 3332 1038
rect 1512 777 1656 807
rect 1209 489 2175 519
rect 129 273 2895 303
rect 1512 201 1656 231
rect 2649 201 3183 231
rect 993 129 1815 159
rect 2433 129 3111 159
rect 417 57 2751 87
rect -20 -30 3332 30
<< metal3 >>
rect 57 360 87 648
rect 129 201 159 303
rect 345 273 375 375
rect 705 360 735 648
rect 417 57 447 231
rect 921 57 951 375
rect 1065 273 1095 375
rect 1209 345 1239 519
rect 1281 273 1311 375
rect 1425 57 1455 375
rect 1785 129 1815 375
rect 1857 201 1887 519
rect 2145 345 2175 519
rect 2361 273 2391 375
rect 2505 57 2535 375
rect 2649 201 2679 375
rect 2721 57 2751 375
rect 2865 273 2895 375
rect 3081 129 3111 375
rect 3153 216 3183 792
use logic_generated_inv_2x  inv0 ~/laygo2_workspace_sky130/magic_layout/logic_generated
timestamp 1704925594
transform 1 0 0 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv1
timestamp 1704925594
transform 1 0 288 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv2
timestamp 1704925594
transform 1 0 1728 0 1 0
box -20 -30 308 1038
use logic_generated_inv_2x  inv3
timestamp 1704925594
transform 1 0 3024 0 1 0
box -20 -30 308 1038
use ntap_fast_boundary  MNT0_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825115
transform 1 0 1440 0 1 0
box 0 0 72 512
use ntap_fast_boundary  MNT0_IBNDR0
timestamp 1655825115
transform 1 0 1656 0 1 0
box 0 0 72 512
use ntap_fast_center_nf2_v2  MNT0_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656694979
transform 1 0 1512 0 1 0
box -36 143 180 342
use via_M1_M2_0  MNT0_IVTAP10 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1584 0 1 216
box -16 -16 16 16
use via_M1_M2_1  MNT0_IVTIETAP10 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 1512 0 1 0
box -16 -16 16 16
use ptap_fast_boundary  MPT0_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825477
transform 1 0 1440 0 -1 1008
box 0 0 84 512
use ptap_fast_boundary  MPT0_IBNDR0
timestamp 1655825477
transform 1 0 1656 0 -1 1008
box 0 0 84 512
use ptap_fast_center_nf2_v2  MPT0_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656699071
transform 1 0 1512 0 -1 1008
box -36 66 180 342
use via_M1_M2_0  MPT0_IVTAP10
timestamp 1647525606
transform 1 0 1584 0 -1 792
box -16 -16 16 16
use via_M1_M2_1  MPT0_IVTIETAP10
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 1512 0 -1 1008
box -16 -16 16 16
use via_M2_M3_0  NoName_1 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 432 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 936 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 2520 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 1440 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_9
timestamp 1647525786
transform 1 0 2736 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_12
timestamp 1647525786
transform 1 0 1800 0 1 144
box -19 -19 19 19
use via_M2_M3_0  NoName_17
timestamp 1647525786
transform 1 0 3096 0 1 144
box -19 -19 19 19
use via_M2_M3_0  NoName_21
timestamp 1647525786
transform 1 0 3168 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_23
timestamp 1647525786
transform 1 0 2664 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_26
timestamp 1647525786
transform 1 0 144 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_28
timestamp 1647525786
transform 1 0 360 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_30
timestamp 1647525786
transform 1 0 1080 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_32
timestamp 1647525786
transform 1 0 2376 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_34
timestamp 1647525786
transform 1 0 1296 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_36
timestamp 1647525786
transform 1 0 2880 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_39
timestamp 1647525786
transform 1 0 1872 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_41
timestamp 1647525786
transform 1 0 2160 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_43
timestamp 1647525786
transform 1 0 1224 0 1 504
box -19 -19 19 19
use logic_generated_tinv_2x  tinv0 ~/laygo2_workspace_sky130/magic_layout/logic_generated
timestamp 1704925691
transform 1 0 576 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_2x  tinv1
timestamp 1704925691
transform 1 0 2016 0 1 0
box -20 -30 596 1038
use logic_generated_tinv_small_1x  tinv_small0 ~/laygo2_workspace_sky130/magic_layout/logic_generated
timestamp 1704925630
transform 1 0 1152 0 1 0
box -20 -30 452 1038
use logic_generated_tinv_small_1x  tinv_small1
timestamp 1704925630
transform 1 0 2592 0 1 0
box -20 -30 452 1038
use via_M2_M3_0  via_M2_M3_0_0
timestamp 1647525786
transform 1 0 1008 0 1 144
box -19 -19 19 19
use via_M2_M3_0  via_M2_M3_0_1
timestamp 1647525786
transform 1 0 1368 0 1 144
box -19 -19 19 19
use via_M2_M3_0  via_M2_M3_0_2
timestamp 1647525786
transform 1 0 2448 0 1 144
box -19 -19 19 19
use via_M2_M3_0  via_M2_M3_0_3
timestamp 1647525786
transform 1 0 2808 0 1 144
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 CLK
port 1 nsew
flabel metal3 720 504 720 504 0 FreeSans 240 90 0 0 I
port 2 nsew
flabel metal3 3168 504 3168 504 0 FreeSans 240 90 0 0 O
port 3 nsew
flabel metal2 1656 1008 1656 1008 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel metal2 1656 0 1656 0 0 FreeSans 480 0 0 0 VSS
port 5 nsew
<< end >>

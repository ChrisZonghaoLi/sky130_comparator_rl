magic
tech sky130A
magscale 1 2
timestamp 1737400462
<< metal1 >>
rect 402 2696 462 3064
rect 690 2696 750 3064
rect 834 2696 894 3064
rect 1122 2696 1182 3064
rect 1266 2696 1326 3064
rect 1554 2696 1614 3064
rect -750 968 -690 1336
rect -462 968 -402 1336
rect -174 402 -114 1336
rect 114 968 174 1336
rect 402 968 462 1336
rect 690 968 750 1336
rect 1266 968 1326 1336
rect 1554 968 1614 1336
rect 1842 968 1902 1336
rect 2130 402 2190 1336
rect 2418 968 2478 1336
rect 2706 968 2766 1336
rect -750 -40 -690 328
rect -462 -40 -402 328
rect 114 -40 174 328
rect 402 -40 462 328
rect 690 -40 750 328
rect 978 -40 1038 328
rect 1266 -40 1326 328
rect 1554 -40 1614 328
rect 1842 -40 1902 328
rect 2418 -40 2478 328
rect 2706 -40 2766 328
<< metal2 >>
rect 228 2964 1788 3084
rect 396 2562 894 2622
rect 1122 2562 1620 2622
rect 396 2274 1620 2334
rect -652 1698 652 1758
rect 1364 1698 2668 1758
rect -652 1410 894 1470
rect 1122 1410 2668 1470
rect -884 1038 884 1068
rect -894 978 884 1038
rect -884 948 884 978
rect 1132 1038 2900 1068
rect 1132 978 2910 1038
rect 1132 948 2900 978
rect 212 690 1804 750
rect -174 402 2190 462
rect -924 -60 2940 60
<< metal3 >>
rect 834 1410 894 2622
rect 978 690 1038 2334
rect 1122 1410 1182 2622
use nmos13_fast_boundary  M1_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 -864 0 1 1008
box 0 0 144 1008
use nmos13_fast_boundary  M1_IBNDR0
timestamp 1655824928
transform 1 0 720 0 1 1008
box 0 0 144 1008
use nfet_01v8_0p84_nf2  M1_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 4 288 0 0 1008
timestamp 1706136540
transform 1 0 -720 0 1 1008
box -92 287 379 721
use via_M1_M2_0  M1_IVD0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 4 288 0 0 1008
timestamp 1709070663
transform 1 0 -576 0 1 1440
box -32 -32 32 32
use via_M1_M2_0  M1_IVG0
array 0 4 288 0 0 1008
timestamp 1709070663
transform 1 0 -576 0 1 1728
box -32 -32 32 32
use via_M1_M2_1  M1_IVTIED0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 5 288 0 0 1008
timestamp 1647525606
transform 1 0 -720 0 1 1008
box -32 -32 32 32
use nmos13_fast_boundary  M2_IBNDL0
timestamp 1655824928
transform 1 0 1152 0 1 1008
box 0 0 144 1008
use nmos13_fast_boundary  M2_IBNDR0
timestamp 1655824928
transform 1 0 2736 0 1 1008
box 0 0 144 1008
use nfet_01v8_0p84_nf2  M2_IM0
array 0 4 288 0 0 1008
timestamp 1706136540
transform 1 0 1296 0 1 1008
box -92 287 379 721
use via_M1_M2_0  M2_IVD0
array 0 4 288 0 0 1008
timestamp 1709070663
transform 1 0 1440 0 1 1440
box -32 -32 32 32
use via_M1_M2_0  M2_IVG0
array 0 4 288 0 0 1008
timestamp 1709070663
transform 1 0 1440 0 1 1728
box -32 -32 32 32
use via_M1_M2_1  M2_IVTIED0
array 0 5 288 0 0 1008
timestamp 1647525606
transform 1 0 1296 0 1 1008
box -32 -32 32 32
use pmos13_fast_boundary  M3_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 288 0 -1 3024
box 0 0 144 1008
use pmos13_fast_boundary  M3_IBNDR0
timestamp 1655825313
transform 1 0 720 0 -1 3024
box 0 0 144 1008
use pfet_01v8_0p42_nf2  M3_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1706648821
transform 1 0 432 0 -1 3024
box -92 132 380 757
use via_M1_M2_0  M3_IVD0
timestamp 1709070663
transform 1 0 576 0 -1 2592
box -32 -32 32 32
use via_M1_M2_0  M3_IVG0
timestamp 1709070663
transform 1 0 576 0 -1 2304
box -32 -32 32 32
use via_M1_M2_1  M3_IVTIED0
array 0 1 288 0 0 -1008
timestamp 1647525606
transform 1 0 432 0 -1 3024
box -32 -32 32 32
use pmos13_fast_boundary  M4_IBNDL0
timestamp 1655825313
transform 1 0 1152 0 -1 3024
box 0 0 144 1008
use pmos13_fast_boundary  M4_IBNDR0
timestamp 1655825313
transform 1 0 1584 0 -1 3024
box 0 0 144 1008
use pfet_01v8_0p42_nf2  M4_IM0
timestamp 1706648821
transform 1 0 1296 0 -1 3024
box -92 132 380 757
use via_M1_M2_0  M4_IVD0
timestamp 1709070663
transform 1 0 1440 0 -1 2592
box -32 -32 32 32
use via_M1_M2_0  M4_IVG0
timestamp 1709070663
transform 1 0 1440 0 -1 2304
box -32 -32 32 32
use via_M1_M2_1  M4_IVTIED0
array 0 1 288 0 0 -1008
timestamp 1647525606
transform 1 0 1296 0 -1 3024
box -32 -32 32 32
use nmos13_fast_boundary  M5_IBNDL0
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 144 1008
use nmos13_fast_boundary  M5_IBNDR0
timestamp 1655824928
transform 1 0 1872 0 1 0
box 0 0 144 1008
use nfet_01v8_0p42_nf2  M5_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 5 288 0 0 1008
timestamp 1706310608
transform 1 0 144 0 1 0
box -92 287 379 757
use via_M1_M2_0  M5_IVD0
array 0 5 288 0 0 1008
timestamp 1709070663
transform 1 0 288 0 1 432
box -32 -32 32 32
use via_M1_M2_0  M5_IVG0
array 0 5 288 0 0 1008
timestamp 1709070663
transform 1 0 288 0 1 720
box -32 -32 32 32
use via_M1_M2_1  M5_IVTIED0
array 0 6 288 0 0 1008
timestamp 1647525606
transform 1 0 144 0 1 0
box -32 -32 32 32
use via_M2_M3_0  NoName_4 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1709070663
transform 1 0 1008 0 1 720
box -38 -38 38 38
use via_M2_M3_0  NoName_6
timestamp 1709070663
transform 1 0 1008 0 1 2304
box -38 -38 38 38
use via_M1_M2_0  NoName_8
timestamp 1709070663
transform 1 0 -144 0 1 432
box -32 -32 32 32
use via_M1_M2_0  NoName_9
timestamp 1709070663
transform 1 0 -144 0 1 1008
box -32 -32 32 32
use via_M1_M2_0  NoName_12
timestamp 1709070663
transform 1 0 2160 0 1 432
box -32 -32 32 32
use via_M1_M2_0  NoName_13
timestamp 1709070663
transform 1 0 2160 0 1 1008
box -32 -32 32 32
use via_M2_M3_0  NoName_17
timestamp 1709070663
transform 1 0 864 0 1 1440
box -38 -38 38 38
use via_M2_M3_0  NoName_18
timestamp 1709070663
transform 1 0 864 0 1 2592
box -38 -38 38 38
use via_M1_M2_0  NoName_20
timestamp 1709070663
transform 1 0 576 0 1 2592
box -32 -32 32 32
use via_M2_M3_0  NoName_23
timestamp 1709070663
transform 1 0 1152 0 1 1440
box -38 -38 38 38
use via_M2_M3_0  NoName_24
timestamp 1709070663
transform 1 0 1152 0 1 2592
box -38 -38 38 38
use via_M1_M2_0  NoName_27
timestamp 1709070663
transform 1 0 1440 0 1 2592
box -32 -32 32 32
use pwell_boundary_0p72_5p04  Ntap_0_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1706900133
transform 1 0 -864 0 1 0
box 0 0 144 1008
use pwell_boundary_0p72_5p04  Ntap_0_IBNDR0
timestamp 1706900133
transform 1 0 -432 0 1 0
box 0 0 144 1008
use ntap_nf2  Ntap_0_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1706909938
transform 1 0 -720 0 1 0
box -72 0 360 1008
use via_M1_M2_1  Ntap_0_IVTIETAP10
array 0 1 288 0 0 1008
timestamp 1647525606
transform 1 0 -720 0 1 0
box -32 -32 32 32
use pwell_boundary_0p72_5p04  Ntap_1_IBNDL0
timestamp 1706900133
transform 1 0 2304 0 1 0
box 0 0 144 1008
use pwell_boundary_0p72_5p04  Ntap_1_IBNDR0
timestamp 1706900133
transform 1 0 2736 0 1 0
box 0 0 144 1008
use ntap_nf2  Ntap_1_IM0
timestamp 1706909938
transform 1 0 2448 0 1 0
box -72 0 360 1008
use via_M1_M2_1  Ntap_1_IVTIETAP10
array 0 1 288 0 0 1008
timestamp 1647525606
transform 1 0 2448 0 1 0
box -32 -32 32 32
use nwell_boundary_0p72_5p04  Nwell_fill_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1706900718
transform 1 0 864 0 -1 3024
box 0 0 168 1008
use nwell_boundary_0p72_5p04  Nwell_fill_IBNDR0
timestamp 1706900718
transform 1 0 1296 0 -1 3024
box 0 0 168 1008
use nwell_1p44_5p04  Nwell_fill_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1706848148
transform 1 0 1008 0 -1 3024
box 0 0 288 1008
use nwell_boundary_0p72_5p04  Nwell_M3_IBNDL0
timestamp 1706900718
transform 1 0 288 0 -1 3024
box 0 0 168 1008
use nwell_boundary_0p72_5p04  Nwell_M3_IBNDR0
timestamp 1706900718
transform 1 0 720 0 -1 3024
box 0 0 168 1008
use nwell_1p44_5p04  Nwell_M3_IM0
timestamp 1706848148
transform 1 0 432 0 -1 3024
box 0 0 288 1008
use nwell_boundary_0p72_5p04  Nwell_M4_IBNDL0
timestamp 1706900718
transform 1 0 1152 0 -1 3024
box 0 0 168 1008
use nwell_boundary_0p72_5p04  Nwell_M4_IBNDR0
timestamp 1706900718
transform 1 0 1584 0 -1 3024
box 0 0 168 1008
use nwell_1p44_5p04  Nwell_M4_IM0
timestamp 1706848148
transform 1 0 1296 0 -1 3024
box 0 0 288 1008
use ptap_nf2  Ptap_0_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1706911696
transform 1 0 864 0 -1 3024
box -72 0 360 1008
use via_M1_M2_1  Ptap_0_IVTIETAP10
array 0 1 288 0 0 -1008
timestamp 1647525606
transform 1 0 864 0 -1 3024
box -32 -32 32 32
use pwell_boundary_0p72_5p04  Pwell_fill1_IBNDL0
timestamp 1706900133
transform 1 0 864 0 1 1008
box 0 0 144 1008
use pwell_boundary_0p72_5p04  Pwell_fill1_IBNDR0
timestamp 1706900133
transform 1 0 1296 0 1 1008
box 0 0 144 1008
use pwell_1p44_5p04  Pwell_fill1_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1706848095
transform 1 0 1008 0 1 1008
box 0 0 288 1008
use pwell_boundary_0p72_5p04  Pwell_fill2_IBNDL0
timestamp 1706900133
transform 1 0 -288 0 1 0
box 0 0 144 1008
use pwell_boundary_0p72_5p04  Pwell_fill2_IBNDR0
timestamp 1706900133
transform 1 0 144 0 1 0
box 0 0 144 1008
use pwell_1p44_5p04  Pwell_fill2_IM0
timestamp 1706848095
transform 1 0 -144 0 1 0
box 0 0 288 1008
use pwell_boundary_0p72_5p04  Pwell_fill3_IBNDL0
timestamp 1706900133
transform 1 0 2016 0 1 0
box 0 0 144 1008
use pwell_boundary_0p72_5p04  Pwell_fill3_IBNDR0
timestamp 1706900133
transform 1 0 2448 0 1 0
box 0 0 144 1008
use pwell_1p44_5p04  Pwell_fill3_IM0
timestamp 1706848095
transform 1 0 2160 0 1 0
box 0 0 288 1008
use pwell_boundary_0p72_5p04  Pwell_M1_IBNDL0
timestamp 1706900133
transform 1 0 -864 0 1 1008
box 0 0 144 1008
use pwell_boundary_0p72_5p04  Pwell_M1_IBNDR0
timestamp 1706900133
transform 1 0 720 0 1 1008
box 0 0 144 1008
use pwell_1p44_5p04  Pwell_M1_IM0
array 0 4 288 0 0 1008
timestamp 1706848095
transform 1 0 -720 0 1 1008
box 0 0 288 1008
use pwell_boundary_0p72_5p04  Pwell_M2_IBNDL0
timestamp 1706900133
transform 1 0 1152 0 1 1008
box 0 0 144 1008
use pwell_boundary_0p72_5p04  Pwell_M2_IBNDR0
timestamp 1706900133
transform 1 0 2736 0 1 1008
box 0 0 144 1008
use pwell_1p44_5p04  Pwell_M2_IM0
array 0 4 288 0 0 1008
timestamp 1706848095
transform 1 0 1296 0 1 1008
box 0 0 288 1008
use pwell_boundary_0p72_5p04  Pwell_M5_IBNDL0
timestamp 1706900133
transform 1 0 0 0 1 0
box 0 0 144 1008
use pwell_boundary_0p72_5p04  Pwell_M5_IBNDR0
timestamp 1706900133
transform 1 0 1872 0 1 0
box 0 0 144 1008
use pwell_1p44_5p04  Pwell_M5_IM0
array 0 5 288 0 0 1008
timestamp 1706848095
transform 1 0 144 0 1 0
box 0 0 288 1008
<< labels >>
flabel metal2 1008 720 1008 720 0 FreeSans 480 0 0 0 CLK
port 1 nsew
flabel metal3 864 2016 864 2016 0 FreeSans 480 90 0 0 Di_n
port 2 nsew
flabel metal3 1152 2016 1152 2016 0 FreeSans 480 90 0 0 Di_p
port 3 nsew
flabel metal2 1008 3024 1008 3024 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel metal2 1008 0 1008 0 0 FreeSans 480 0 0 0 VSS
port 5 nsew
flabel metal2 2016 1728 2016 1728 0 FreeSans 480 0 0 0 Vin_n
port 6 nsew
flabel metal2 0 1728 0 1728 0 FreeSans 480 0 0 0 Vin_p
port 7 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1706136540
<< pwell >>
rect -92 401 379 641
<< nmos >>
rect 57 437 87 605
rect 200 437 230 605
<< ndiff >>
rect -56 583 57 605
rect -56 543 -20 583
rect 20 543 57 583
rect -56 499 57 543
rect -56 459 -20 499
rect 20 459 57 499
rect -56 437 57 459
rect 87 583 200 605
rect 87 543 124 583
rect 164 543 200 583
rect 87 499 200 543
rect 87 459 124 499
rect 164 459 200 499
rect 87 437 200 459
rect 230 583 343 605
rect 230 543 268 583
rect 308 543 343 583
rect 230 499 343 543
rect 230 459 268 499
rect 308 459 343 499
rect 230 437 343 459
<< ndiffc >>
rect -20 543 20 583
rect -20 459 20 499
rect 124 543 164 583
rect 124 459 164 499
rect 268 543 308 583
rect 268 459 308 499
<< poly >>
rect 57 701 230 721
rect 57 661 77 701
rect 117 661 170 701
rect 210 661 230 701
rect 57 641 230 661
rect 57 605 87 641
rect 200 605 230 641
rect 57 401 87 437
rect 200 401 230 437
<< polycont >>
rect 77 661 117 701
rect 170 661 210 701
<< locali >>
rect 57 701 230 721
rect 57 661 77 701
rect 117 661 170 701
rect 210 661 230 701
rect 57 641 230 661
rect -30 583 30 599
rect -30 543 -20 583
rect 20 543 30 583
rect -30 499 30 543
rect -30 459 -20 499
rect 20 459 30 499
rect -30 443 30 459
rect 114 583 174 599
rect 114 543 124 583
rect 164 543 174 583
rect 114 499 174 543
rect 114 459 124 499
rect 164 459 174 499
rect 114 443 174 459
rect 258 583 318 599
rect 258 543 268 583
rect 308 543 318 583
rect 258 499 318 543
rect 258 459 268 499
rect 308 459 318 499
rect 258 443 318 459
<< viali >>
rect 77 661 117 701
rect 170 661 210 701
rect -20 543 20 583
rect -20 459 20 499
rect 124 543 164 583
rect 124 459 164 499
rect 268 543 308 583
rect 268 459 308 499
<< metal1 >>
rect 57 701 230 721
rect 57 661 77 701
rect 117 661 170 701
rect 210 661 230 701
rect 57 641 230 661
rect -30 583 30 599
rect -30 543 -20 583
rect 20 543 30 583
rect -30 499 30 543
rect -30 459 -20 499
rect 20 459 30 499
rect -30 287 30 459
rect 114 583 174 599
rect 114 543 124 583
rect 164 543 174 583
rect 114 499 174 543
rect 114 459 124 499
rect 164 459 174 499
rect 114 287 174 459
rect 258 583 318 599
rect 258 543 268 583
rect 308 543 318 583
rect 258 499 318 543
rect 258 459 268 499
rect 308 459 318 499
rect 258 287 318 459
<< end >>

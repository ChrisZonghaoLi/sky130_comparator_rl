magic
tech sky130A
timestamp 1706900133
<< pwell >>
rect 0 0 72 504
<< end >>

magic
tech sky130A
timestamp 1705618273
<< checkpaint >>
rect -650 -660 1370 1668
<< metal1 >>
rect 57 844 87 1028
rect 201 844 231 1028
rect 345 844 375 1028
rect 489 844 519 1028
rect 633 844 663 1028
rect 57 -20 87 164
rect 201 -20 231 164
rect 345 -20 375 164
rect 489 -20 519 164
rect 633 -20 663 164
<< metal2 >>
rect -20 978 740 1038
rect 106 777 614 807
rect 62 633 614 663
rect 62 345 614 375
rect 106 201 614 231
rect -20 -30 740 30
<< metal3 >>
rect 57 345 87 663
rect 561 201 591 807
use nmos13_fast_boundary  MN0_IBNDL0 /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655824928
transform 1 0 0 0 1 0
box 0 0 72 504
use nmos13_fast_boundary  MN0_IBNDR0
timestamp 1655824928
transform 1 0 648 0 1 0
box 0 0 72 504
use nmos13_fast_center_nf2  MN0_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 3 144 0 0 504
timestamp 1654175211
transform 1 0 72 0 1 0
box -46 143 190 378
use via_M1_M2_0  MN0_IVD0 /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 3 144 0 0 504
timestamp 1647525606
transform 1 0 144 0 1 216
box -16 -16 16 16
use via_M1_M2_0  MN0_IVG0
array 0 3 144 0 0 504
timestamp 1647525606
transform 1 0 144 0 1 360
box -16 -16 16 16
use via_M1_M2_1  MN0_IVTIED0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 4 144 0 0 504
timestamp 1647525606
transform 1 0 72 0 1 0
box -16 -16 16 16
use pmos13_fast_boundary  MP0_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825313
transform 1 0 0 0 -1 1008
box 0 0 72 504
use pmos13_fast_boundary  MP0_IBNDR0
timestamp 1655825313
transform 1 0 648 0 -1 1008
box 0 0 72 504
use pmos13_fast_center_nf2  MP0_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 3 144 0 0 -504
timestamp 1654091791
transform 1 0 72 0 -1 1008
box -46 66 190 378
use via_M1_M2_0  MP0_IVD0
array 0 3 144 0 0 -504
timestamp 1647525606
transform 1 0 144 0 -1 792
box -16 -16 16 16
use via_M1_M2_0  MP0_IVG0
array 0 3 144 0 0 -504
timestamp 1647525606
transform 1 0 144 0 -1 648
box -16 -16 16 16
use via_M1_M2_1  MP0_IVTIED0
array 0 4 144 0 0 -504
timestamp 1647525606
transform 1 0 72 0 -1 1008
box -16 -16 16 16
use via_M2_M3_0  NoName_1 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 72 0 1 360
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 72 0 1 648
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 576 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 576 0 1 792
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 I
port 1 nsew
flabel metal3 576 504 576 504 0 FreeSans 240 90 0 0 O
port 2 nsew
flabel metal2 360 1008 360 1008 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal2 360 0 360 0 0 FreeSans 480 0 0 0 VSS
port 4 nsew
<< end >>

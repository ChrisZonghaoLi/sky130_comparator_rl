* NGSPICE file created from comparator_flat.ext - technology: sky130A

.subckt comparator_flat CLK VDD VSS Vin_p Vin_n Di_p Di_n Vout_n CLK_bar Vout_p
X0 VDD CLK_bar latch.inv1.VDD VDD sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X1 Vout_p Vout_n latch.inv1.VDD VDD sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X2 Di_n Vin_p a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X3 latch.inv1.VDD CLK_bar VDD VDD sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X4 a_88_n1613# Vin_p Di_n VSS sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X5 VDD CLK_bar latch.inv1.VDD VDD sky130_fd_pr__pfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X6 Vout_p Di_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X7 a_88_n1613# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X8 a_88_n1613# Vin_p Di_n VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X9 a_88_n1613# Vin_n Di_p VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X10 VSS CLK a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X11 Di_p Vin_n a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X12 Di_p CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X13 a_88_n1613# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X14 VDD CLK Di_p VDD sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X15 a_88_n1613# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X16 VSS CLK a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X17 a_88_n1613# Vin_p Di_n VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X18 latch.inv1.VDD Vout_p Vout_n VDD sky130_fd_pr__pfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X19 Di_n CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X20 Vout_n Vout_p VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X21 VSS Di_n Vout_p VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X22 Di_p Vin_n a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X23 VDD CLK Di_n VDD sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X24 a_88_n1613# Vin_n Di_p VSS sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X25 latch.inv1.VDD CLK_bar VDD VDD sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X26 VSS CLK a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X27 Di_n Vin_p a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X28 Di_n Vin_p a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X29 Vout_n Di_p VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X30 a_88_n1613# Vin_p Di_n VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X31 a_88_n1613# Vin_p Di_n VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X32 a_88_n1613# Vin_n Di_p VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X33 a_88_n1613# Vin_n Di_p VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X34 Di_n Vin_p a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X35 Di_p Vin_n a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X36 latch.inv1.VDD CLK_bar VDD VDD sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X37 latch.inv1.VDD Vout_n Vout_p VDD sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X38 VSS Vout_p Vout_n VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X39 Di_p Vin_n a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X40 VDD CLK_bar latch.inv1.VDD VDD sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X41 Vout_n Vout_p latch.inv1.VDD VDD sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X42 latch.inv1.VDD Vout_p Vout_n VDD sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X43 a_88_n1613# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X44 a_88_n1613# Vin_p Di_n VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X45 VSS Di_p Vout_n VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X46 VSS CLK a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X47 latch.inv1.VDD Vout_n Vout_p VDD sky130_fd_pr__pfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X48 Vout_p Vout_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X49 a_88_n1613# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X50 Vout_n Vout_p latch.inv1.VDD VDD sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X51 VSS CLK a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X52 Di_p Vin_n a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X53 Di_n Vin_p a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X54 a_88_n1613# Vin_n Di_p VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X55 Vout_p Vout_n latch.inv1.VDD VDD sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X56 Di_n Vin_p a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X57 a_88_n1613# Vin_n Di_p VSS sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X58 VSS Vout_n Vout_p VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X59 Di_p Vin_n a_88_n1613# VSS sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
.ends


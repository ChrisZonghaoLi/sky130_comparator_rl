magic
tech sky130A
magscale 1 2
timestamp 1706306204
<< nwell >>
rect -92 383 236 551
<< pmos >>
rect 57 425 87 509
<< pdiff >>
rect -56 487 57 509
rect -56 447 -20 487
rect 20 447 57 487
rect -56 425 57 447
rect 87 487 200 509
rect 87 447 124 487
rect 164 447 200 487
rect 87 425 200 447
<< pdiffc >>
rect -20 447 20 487
rect 124 447 164 487
<< poly >>
rect 32 605 112 625
rect 32 565 52 605
rect 92 565 112 605
rect 32 545 112 565
rect 57 509 87 545
rect 57 389 87 425
<< polycont >>
rect 52 565 92 605
<< locali >>
rect 32 605 112 625
rect 32 565 52 605
rect 92 565 112 605
rect 32 545 112 565
rect -30 487 30 503
rect -30 447 -20 487
rect 20 447 30 487
rect -30 431 30 447
rect 114 487 174 503
rect 114 447 124 487
rect 164 447 174 487
rect 114 431 174 447
<< viali >>
rect 52 565 92 605
rect -20 447 20 487
rect 124 447 164 487
<< metal1 >>
rect 32 605 112 625
rect 32 565 52 605
rect 92 565 112 605
rect 32 545 112 565
rect -30 487 30 503
rect -30 447 -20 487
rect 20 447 30 487
rect -30 383 30 447
rect 114 487 174 503
rect 114 447 124 487
rect 164 447 174 487
rect 114 383 174 447
<< end >>

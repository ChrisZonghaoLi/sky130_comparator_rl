.param W_M1=8.189754198193551
.param W_M3=0.6693031996488568
.param W_M5=4.729764678701758
.param W_M6=1.0326698946952817
.param W_M7=0.5163349473476408
.param W_M10=0.752667883634567
.param W_M12=9.594074639081956
.param W_M2=W_M1
.param W_M4=W_M3
.param W_M9=W_M6
.param W_M8=W_M7
.param W_M11=W_M10
.param Vcm=0.9008961886167527
.param VDD=1.8
.param Vin=0.05
.param Vin_min=0.0001
.param CL=2e-14
.param Tclk=1e-09
.param Tclk_pk=4.5e-10
.param Tdelay=2e-10
.param Tdelay_bar=7.000000000000001e-10
.param Tr=5.000000000000001e-11
.param Tf=5.000000000000001e-11

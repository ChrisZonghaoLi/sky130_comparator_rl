magic
tech sky130A
timestamp 1704925973
<< checkpaint >>
rect -650 -660 5114 1668
<< metal1 >>
rect 2073 844 2103 1028
rect 2217 844 2247 1028
rect 2073 -20 2103 164
rect 2217 -20 2247 164
<< metal2 >>
rect -20 978 4484 1038
rect 2088 777 2232 807
rect 1785 489 2895 519
rect 273 273 3903 303
rect 2088 201 2232 231
rect 3657 201 4335 231
rect 1569 129 2391 159
rect 3441 129 4119 159
rect 705 57 3759 87
rect -20 -30 4484 30
<< metal3 >>
rect 57 360 87 648
rect 273 201 303 303
rect 489 273 519 375
rect 993 360 1023 648
rect 705 57 735 231
rect 1497 57 1527 375
rect 1641 273 1671 375
rect 1785 345 1815 519
rect 1857 273 1887 375
rect 2001 57 2031 375
rect 2361 129 2391 375
rect 2577 201 2607 519
rect 2865 345 2895 519
rect 3369 273 3399 375
rect 3513 57 3543 375
rect 3657 201 3687 375
rect 3729 57 3759 375
rect 3873 273 3903 375
rect 4089 129 4119 375
rect 4305 216 4335 792
use logic_generated_inv_4x  inv0 ~/laygo2_workspace_sky130/magic_layout/logic_generated
timestamp 1704925594
transform 1 0 0 0 1 0
box -20 -30 452 1038
use logic_generated_inv_4x  inv1
timestamp 1704925594
transform 1 0 432 0 1 0
box -20 -30 452 1038
use logic_generated_inv_4x  inv2
timestamp 1704925594
transform 1 0 2304 0 1 0
box -20 -30 452 1038
use logic_generated_inv_4x  inv3
timestamp 1704925594
transform 1 0 4032 0 1 0
box -20 -30 452 1038
use ntap_fast_boundary  MNT0_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825115
transform 1 0 2016 0 1 0
box 0 0 72 512
use ntap_fast_boundary  MNT0_IBNDR0
timestamp 1655825115
transform 1 0 2232 0 1 0
box 0 0 72 512
use ntap_fast_center_nf2_v2  MNT0_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656694979
transform 1 0 2088 0 1 0
box -36 143 180 342
use via_M1_M2_0  MNT0_IVTAP10 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 2160 0 1 216
box -16 -16 16 16
use via_M1_M2_1  MNT0_IVTIETAP10 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
array 0 1 144 0 0 504
timestamp 1647525606
transform 1 0 2088 0 1 0
box -16 -16 16 16
use ptap_fast_boundary  MPT0_IBNDL0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1655825477
transform 1 0 2016 0 -1 1008
box 0 0 84 512
use ptap_fast_boundary  MPT0_IBNDR0
timestamp 1655825477
transform 1 0 2232 0 -1 1008
box 0 0 84 512
use ptap_fast_center_nf2_v2  MPT0_IM0 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1656699071
transform 1 0 2088 0 -1 1008
box -36 66 180 342
use via_M1_M2_0  MPT0_IVTAP10
timestamp 1647525606
transform 1 0 2160 0 -1 792
box -16 -16 16 16
use via_M1_M2_1  MPT0_IVTIETAP10
array 0 1 144 0 0 -504
timestamp 1647525606
transform 1 0 2088 0 -1 1008
box -16 -16 16 16
use via_M2_M3_0  NoName_1 ~/laygo2_workspace_sky130/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 720 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_3
timestamp 1647525786
transform 1 0 1512 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_5
timestamp 1647525786
transform 1 0 3528 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_7
timestamp 1647525786
transform 1 0 2016 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_9
timestamp 1647525786
transform 1 0 3744 0 1 72
box -19 -19 19 19
use via_M2_M3_0  NoName_12
timestamp 1647525786
transform 1 0 2376 0 1 144
box -19 -19 19 19
use via_M2_M3_0  NoName_17
timestamp 1647525786
transform 1 0 4104 0 1 144
box -19 -19 19 19
use via_M2_M3_0  NoName_19
timestamp 1647525786
transform 1 0 3816 0 1 144
box -19 -19 19 19
use via_M2_M3_0  NoName_23
timestamp 1647525786
transform 1 0 3672 0 1 216
box -19 -19 19 19
use via_M2_M3_0  NoName_26
timestamp 1647525786
transform 1 0 288 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_28
timestamp 1647525786
transform 1 0 504 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_30
timestamp 1647525786
transform 1 0 1656 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_32
timestamp 1647525786
transform 1 0 3384 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_34
timestamp 1647525786
transform 1 0 1872 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_36
timestamp 1647525786
transform 1 0 3888 0 1 288
box -19 -19 19 19
use via_M2_M3_0  NoName_39
timestamp 1647525786
transform 1 0 2592 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_41
timestamp 1647525786
transform 1 0 2880 0 1 504
box -19 -19 19 19
use via_M2_M3_0  NoName_43
timestamp 1647525786
transform 1 0 1800 0 1 504
box -19 -19 19 19
use logic_generated_tinv_4x  tinv0 ~/laygo2_workspace_sky130/magic_layout/logic_generated
timestamp 1704925691
transform 1 0 864 0 1 0
box -20 -30 884 1038
use logic_generated_tinv_4x  tinv1
timestamp 1704925691
transform 1 0 2736 0 1 0
box -20 -30 884 1038
use logic_generated_tinv_small_1x  tinv_small0 ~/laygo2_workspace_sky130/magic_layout/logic_generated
timestamp 1704925630
transform 1 0 1728 0 1 0
box -20 -30 452 1038
use logic_generated_tinv_small_1x  tinv_small1
timestamp 1704925630
transform 1 0 3600 0 1 0
box -20 -30 452 1038
use via_M2_M3_0  via_M2_M3_0_0
timestamp 1647525786
transform 1 0 1584 0 1 144
box -19 -19 19 19
use via_M2_M3_0  via_M2_M3_0_1
timestamp 1647525786
transform 1 0 1944 0 1 144
box -19 -19 19 19
use via_M2_M3_0  via_M2_M3_0_2
timestamp 1647525786
transform 1 0 3456 0 1 144
box -19 -19 19 19
use via_M2_M3_0  via_M2_M3_0_3
timestamp 1647525786
transform 1 0 4320 0 1 216
box -19 -19 19 19
<< labels >>
flabel metal3 72 504 72 504 0 FreeSans 240 90 0 0 CLK
port 1 nsew
flabel metal3 1008 504 1008 504 0 FreeSans 240 90 0 0 I
port 2 nsew
flabel metal3 4320 504 4320 504 0 FreeSans 240 90 0 0 O
port 3 nsew
flabel metal2 2232 1008 2232 1008 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel metal2 2232 0 2232 0 0 FreeSans 480 0 0 0 VSS
port 5 nsew
<< end >>

.param W_M1=8.4
.param W_M3=0.84
.param W_M5=5.04
.param W_M6=1.68
.param W_M7=0.84
.param W_M10=0.84
.param W_M12=10.08
.param W_M2=W_M1
.param W_M4=W_M3
.param W_M9=W_M6
.param W_M8=W_M7
.param W_M11=W_M10
.param Vcm=0.91
.param VDD=1.8
.param Vin=0.05
.param Vin_min=0.0001
.param CL=2e-14
.param Tclk=1e-09
.param Tclk_pk=4.5e-10
.param Tdelay=2e-10
.param Tdelay_bar=7.000000000000001e-10
.param Tr=5.000000000000001e-11
.param Tf=5.000000000000001e-11

.param W_M1=9.52179530620575
.param W_M3=0.8479869997501375
.param W_M5=9.94891750752926
.param W_M6=0.5590121358633038
.param W_M7=0.6923666799068453
.param W_M10=1.5256951802968977
.param W_M12=6.560755328834057
.param W_M2=W_M1
.param W_M4=W_M3
.param W_M9=W_M6
.param W_M8=W_M7
.param W_M11=W_M10
.param Vcm=0.9030247986316682
.param VDD=1.8
.param Vin=0.05
.param Vin_min=0.0001
.param CL=2e-14
.param Tclk=1e-09
.param Tclk_pk=4.5e-10
.param Tdelay=2e-10
.param Tdelay_bar=7.000000000000001e-10
.param Tr=5.000000000000001e-11
.param Tf=5.000000000000001e-11


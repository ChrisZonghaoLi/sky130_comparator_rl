.param W_M1=1.0
.param W_M3=1.0
.param W_M5=1.0
.param W_M7=1.0
.param W_M8=1.0
.param W_M10=1.0
.param W_M2=W_M1
.param W_M4=W_M3
.param W_M6=W_M5
.param W_M9=W_M8
.param W_M11=W_M10
.param Vcm=1.1
.param VDD=1.8
.param Vin=0.05
.param Vin_min=0.0001
.param CL=2e-14
.param Tclk=1e-09
.param Tclk_pk=4.5e-10
.param Tdelay=2e-10
.param Tr=5.000000000000001e-11
.param Tf=5.000000000000001e-11


** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp_pex_tb.sch
**.subckt double_tail_comp_pex_tb Di_n Di_p Vout_n Vout_p Q Q_bar Di_n_mc Di_p_mc Vout_n_mc
*+ Vout_p_mc Di_n_ms Di_p_ms Vout_n_ms Vout_p_ms Di_n_kn Di_p_kn Vout_n_kn Vout_p_kn
*.opin Di_n
*.opin Di_p
*.opin Vout_n
*.opin Vout_p
*.opin Q
*.opin Q_bar
*.opin Di_n_mc
*.opin Di_p_mc
*.opin Vout_n_mc
*.opin Vout_p_mc
*.opin Di_n_ms
*.opin Di_p_ms
*.opin Vout_n_ms
*.opin Vout_p_ms
*.opin Di_n_kn
*.opin Di_p_kn
*.opin Vout_n_kn
*.opin Vout_p_kn
x1 net1 Vclk_bar Vout_n Vout_p Di_n Di_p Vcm net10 Vclk GND double_tail_comp
VDD net1 net9 VDD
Vclk Vclk GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar Vclk_bar GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm Vcm GND dc Vcm
Vdiff net10 Vcm dc Vin
C2 Q_bar GND 10f m=1
C3 Q GND 10f m=1
x2 net17 Vout_n Q Vout_p Q_bar RS_latch
x3 net4 net3 Vout_n_mc Vout_p_mc Di_n_mc Di_p_mc net2 Vsc net15 GND double_tail_comp
VDD2 net4 GND VDD
Vclk2 net15 GND PULSE(0 VDD 0 Tr Tf Tclk_pk Tclk 0)
Vclk_bar2 net3 GND PULSE(0 VDD Tclk_pk Tr Tf Tclk_pk Tclk 0)
Vcm2 net2 GND dc Vcm
ASRC1 %v([ Vsc ]) filesrc
x4 net8 net7 Vout_n_ms Vout_p_ms Di_n_ms Di_p_ms net5 net6 net16 GND double_tail_comp
VDD3 net8 GND VDD
Vclk3 net16 GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar3 net7 GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm3 net5 GND dc Vcm
Vdiff2 net6 net5 dc Vin_min
VDD_latch net17 GND VDD
Rdummy net9 GND 1 m=1
x5 net13 net12 Vout_n_kn Vout_p_kn Di_n_kn Di_p_kn Vn_kn Vp_kn net18 GND double_tail_comp
VDD4 net13 GND VDD
Vclk4 net18 GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar5 net12 GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm4 net11 GND dc Vcm
Vdiff4 net14 net11 dc Vin
Rdummyn net11 Vn_kn 8k m=1
Rdummyp net14 Vp_kn 8k m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



*.OPTIONS maxord=1
*.OPTIONS itl1=200
*.OPTIONS itl2=200
*.OPTIONS itl4=200

* save all voltage and current
.save all
.options savecurrents
.options seed=random

.control
set filetype=ascii
set units=degrees

* RC extracted comparator netlist
.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/sky130_comparator/netgen/double_tail/TCL/double_tail_comparator_pex.spice
* analyses
.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/sky130_comparator/comparator_transfer_learning/pex/simulations/double_tail_comp_pex_tb_analyses.spice
* stimulus variables
.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/sky130_comparator/comparator_transfer_learning/pex/simulations/double_tail_comp_pex_tb_vars.spice

.endc


**** end user architecture code
**.ends

* expanding   symbol:  double_tail_comp.sym # of pins=10
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp.sch
.subckt double_tail_comp VDD CLK_bar Vout_n Vout_p Di_p Di_n Vin_n Vin_p CLK VSS
+ Vout_p
X0 VSS.t36 CLK.t0 a_88_n1613.t11 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X1 a_88_n1613.t7 CLK.t1 VSS.t34 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X2 a_88_n1613.t12 CLK.t2 VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X3 Vout_p.t3 Di_n.t12 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X4 Vout_p.t2 Di_n.t13 VSS.t38 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X5 a_88_n1613.t3 Vin_p.t0 Di_n.t2 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X6 a_88_n1613.t28 Vin_n.t0 Di_p.t11 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X7 Vout_p.t6 Vout_n.t8 VSS.t49 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X8 a_88_n1613.t9 CLK.t3 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X9 Di_p.t10 Vin_n.t1 a_88_n1613.t20 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X10 VSS.t11 Vout_p.t8 Vout_n.t3 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X11 VDD.t34 CLK_bar.t0 latch.inv0.VDD VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X12 a_88_n1613.t5 CLK.t4 VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X13 latch.inv0.VDD Vout_p.t9 Vout_n.t1 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X14 a_88_n1613.t21 Vin_p.t1 Di_n.t7 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X15 VDD.t32 CLK_bar.t1 latch.inv0.VDD VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X16 VSS.t9 Di_n.t14 Vout_p.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X17 Di_p.t9 Vin_n.t2 a_88_n1613.t2 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X18 latch.inv0.VDD CLK_bar.t2 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X19 latch.inv0.VDD CLK_bar.t3 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X20 VSS.t26 CLK.t5 a_88_n1613.t13 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X21 VSS.t53 Di_n.t15 Vout_p.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X22 Di_p.t8 Vin_n.t3 a_88_n1613.t23 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X23 VDD.t11 CLK.t6 Di_p.t0 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X24 latch.inv0.VDD CLK_bar.t4 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X25 VSS.t24 CLK.t7 a_88_n1613.t16 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X26 a_88_n1613.t10 CLK.t8 VSS.t22 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X27 Di_n.t9 Vin_p.t2 a_88_n1613.t26 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X28 Di_n.t6 Vin_p.t3 a_88_n1613.t18 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X29 VSS.t21 CLK.t9 a_88_n1613.t14 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X30 a_88_n1613.t0 Vin_p.t4 Di_n.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X31 a_88_n1613.t1 Vin_p.t5 Di_n.t1 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X32 a_88_n1613.t31 Vin_n.t4 Di_p.t7 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X33 a_88_n1613.t4 Vin_n.t5 Di_p.t6 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X34 latch.inv0.VDD CLK_bar.t5 VDD.t24 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X35 a_88_n1613.t8 CLK.t10 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X36 Di_n.t8 Vin_p.t6 a_88_n1613.t24 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X37 VSS.t54 Vout_n.t9 Vout_p.t7 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X38 Di_p.t5 Vin_n.t6 a_88_n1613.t22 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X39 VSS.t17 CLK.t11 a_88_n1613.t15 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X40 Di_p.t1 CLK.t12 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X41 VDD.t23 CLK_bar.t6 latch.inv0.VDD VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X42 a_88_n1613.t17 Vin_p.t7 Di_n.t5 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X43 Vout_n.t0 Vout_p.t10 latch.inv0.VDD VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X44 VSS.t14 Di_p.t12 Vout_n.t7 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X45 VDD.t21 CLK_bar.t7 latch.inv0.VDD VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X46 Vout_n.t2 Vout_p.t11 VSS.t40 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X47 latch.inv0.VDD CLK_bar.t8 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X48 latch.inv0.VDD Vout_n.t10 Vout_p.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X49 Vout_n.t6 Di_p.t13 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X50 Vout_n.t5 Di_p.t14 VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X51 Di_n.t4 CLK.t13 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X52 VDD.t17 CLK_bar.t9 latch.inv0.VDD VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X53 VDD.t5 CLK.t14 Di_n.t3 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X54 latch.inv0.VDD CLK_bar.t10 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X55 Di_p.t4 Vin_n.t7 a_88_n1613.t29 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X56 VDD.t13 CLK_bar.t11 latch.inv0.VDD VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X57 Di_n.t11 Vin_p.t8 a_88_n1613.t30 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X58 a_88_n1613.t19 Vin_n.t8 Di_p.t3 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X59 Vout_p.t5 Vout_n.t11 latch.inv0.VDD VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X60 VSS.t47 Di_p.t15 Vout_n.t4 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X61 VSS.t15 CLK.t15 a_88_n1613.t6 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X62 Di_n.t10 Vin_p.t9 a_88_n1613.t27 VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X63 a_88_n1613.t25 Vin_n.t9 Di_p.t2 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
R0 CLK.n6 CLK.t13 164.137
R1 CLK.n6 CLK.t14 164.137
R2 CLK.n5 CLK.t12 164.137
R3 CLK.n5 CLK.t6 164.137
R4 CLK.n11 CLK.t0 164.137
R5 CLK.n11 CLK.t4 164.137
R6 CLK.n9 CLK.t15 164.137
R7 CLK.n9 CLK.t3 164.137
R8 CLK.n8 CLK.t11 164.137
R9 CLK.n8 CLK.t2 164.137
R10 CLK.n3 CLK.t7 164.137
R11 CLK.n3 CLK.t1 164.137
R12 CLK.n1 CLK.t9 164.137
R13 CLK.n1 CLK.t8 164.137
R14 CLK.n0 CLK.t5 164.137
R15 CLK.n0 CLK.t10 164.137
R16 CLK.n7 CLK.n6 74.2428
R17 CLK.n7 CLK.n5 74.2428
R18 CLK.n10 CLK.n8 73.9553
R19 CLK.n2 CLK.n0 73.9553
R20 CLK.n12 CLK.n11 73.3637
R21 CLK.n10 CLK.n9 73.3637
R22 CLK.n4 CLK.n3 73.3637
R23 CLK.n2 CLK.n1 73.3637
R24 CLK CLK.n7 8.04877
R25 CLK.n12 CLK.n10 0.592167
R26 CLK.n4 CLK.n2 0.592167
R27 CLK CLK.n12 0.279667
R28 CLK CLK.n4 0.279667
R29 a_88_n1613.n1 a_88_n1613.n16 198.894
R30 a_88_n1613.n1 a_88_n1613.n15 198.894
R31 a_88_n1613.n1 a_88_n1613.n14 198.894
R32 a_88_n1613.n1 a_88_n1613.n13 198.894
R33 a_88_n1613.n0 a_88_n1613.n12 198.894
R34 a_88_n1613.n0 a_88_n1613.n11 198.894
R35 a_88_n1613.n3 a_88_n1613.t4 144.418
R36 a_88_n1613.n2 a_88_n1613.t1 144.418
R37 a_88_n1613.n3 a_88_n1613.t2 143.703
R38 a_88_n1613.n2 a_88_n1613.t26 143.703
R39 a_88_n1613.t27 a_88_n1613.n2 102.689
R40 a_88_n1613.n3 a_88_n1613.n8 102.689
R41 a_88_n1613.n3 a_88_n1613.n9 102.689
R42 a_88_n1613.n3 a_88_n1613.n7 102.689
R43 a_88_n1613.n2 a_88_n1613.n5 102.689
R44 a_88_n1613.n2 a_88_n1613.n4 102.689
R45 a_88_n1613.n10 a_88_n1613.n6 98.1895
R46 a_88_n1613.n18 a_88_n1613.n17 98.1895
R47 a_88_n1613.n16 a_88_n1613.t12 81.4291
R48 a_88_n1613.n15 a_88_n1613.t9 81.4291
R49 a_88_n1613.n14 a_88_n1613.t5 81.4291
R50 a_88_n1613.n13 a_88_n1613.t7 81.4291
R51 a_88_n1613.n12 a_88_n1613.t10 81.4291
R52 a_88_n1613.n11 a_88_n1613.t8 81.4291
R53 a_88_n1613.n16 a_88_n1613.t15 80.0005
R54 a_88_n1613.n15 a_88_n1613.t6 80.0005
R55 a_88_n1613.n14 a_88_n1613.t11 80.0005
R56 a_88_n1613.n13 a_88_n1613.t16 80.0005
R57 a_88_n1613.n12 a_88_n1613.t14 80.0005
R58 a_88_n1613.n11 a_88_n1613.t13 80.0005
R59 a_88_n1613.n8 a_88_n1613.t28 41.4291
R60 a_88_n1613.n9 a_88_n1613.t19 41.4291
R61 a_88_n1613.n7 a_88_n1613.t25 41.4291
R62 a_88_n1613.n6 a_88_n1613.t31 41.4291
R63 a_88_n1613.n17 a_88_n1613.t3 41.4291
R64 a_88_n1613.n5 a_88_n1613.t17 41.4291
R65 a_88_n1613.n4 a_88_n1613.t21 41.4291
R66 a_88_n1613.t0 a_88_n1613.t27 41.4291
R67 a_88_n1613.n8 a_88_n1613.t29 40.7148
R68 a_88_n1613.n9 a_88_n1613.t20 40.7148
R69 a_88_n1613.n7 a_88_n1613.t23 40.7148
R70 a_88_n1613.n6 a_88_n1613.t22 40.7148
R71 a_88_n1613.n17 a_88_n1613.t24 40.7148
R72 a_88_n1613.n5 a_88_n1613.t30 40.7148
R73 a_88_n1613.n4 a_88_n1613.t18 40.7148
R74 a_88_n1613.n0 a_88_n1613.n10 6.58383
R75 a_88_n1613.n18 a_88_n1613.n1 6.58383
R76 a_88_n1613.n10 a_88_n1613.n3 5.4005
R77 a_88_n1613.n2 a_88_n1613.n18 5.4005
R78 a_88_n1613.n1 a_88_n1613.n0 2.95883
R79 VSS.n66 VSS.n17 87233.1
R80 VSS.n65 VSS.n49 37625.4
R81 VSS.n60 VSS.n59 669.847
R82 VSS.n42 VSS.n41 669.847
R83 VSS.n57 VSS.n56 585
R84 VSS.n58 VSS.n57 585
R85 VSS.n16 VSS.n15 585
R86 VSS.n64 VSS.n16 585
R87 VSS.n69 VSS.n68 585
R88 VSS.n68 VSS.n67 585
R89 VSS.n47 VSS.n46 585
R90 VSS.n48 VSS.n47 585
R91 VSS.n20 VSS.n19 585
R92 VSS.n63 VSS.n62 585
R93 VSS.n64 VSS.n63 585
R94 VSS.n61 VSS.n50 585
R95 VSS.n26 VSS.n25 585
R96 VSS.n25 VSS.n24 585
R97 VSS.n23 VSS.n18 585
R98 VSS.n48 VSS.n18 585
R99 VSS.n39 VSS.n38 585
R100 VSS.n40 VSS.n39 585
R101 VSS.n41 VSS.n40 300.947
R102 VSS.n59 VSS.n58 300.947
R103 VSS.n76 VSS.t53 282.651
R104 VSS.n11 VSS.t49 282.651
R105 VSS.n0 VSS.t11 282.651
R106 VSS.n30 VSS.t26 282.651
R107 VSS.n33 VSS.t14 282.651
R108 VSS.n72 VSS.t7 281.223
R109 VSS.n75 VSS.t32 281.223
R110 VSS.n9 VSS.t54 281.223
R111 VSS.n2 VSS.t40 281.223
R112 VSS.n29 VSS.t5 281.223
R113 VSS.t18 VSS.t20 210.98
R114 VSS.t33 VSS.t35 210.98
R115 VSS.t29 VSS.t16 210.98
R116 VSS.t55 VSS.t45 208.07
R117 VSS.t13 VSS.t42 208.07
R118 VSS.t58 VSS.t44 208.07
R119 VSS.t46 VSS.t4 208.07
R120 VSS.t25 VSS.t18 208.07
R121 VSS.t20 VSS.t2 208.07
R122 VSS.t10 VSS.t39 208.07
R123 VSS.t23 VSS.t33 208.07
R124 VSS.t35 VSS.t27 208.07
R125 VSS.t27 VSS.t48 208.07
R126 VSS.t1 VSS.t29 208.07
R127 VSS.t16 VSS.t31 208.07
R128 VSS.t52 VSS.t37 208.07
R129 VSS.t41 VSS.t51 208.07
R130 VSS.t8 VSS.t6 208.07
R131 VSS.t3 VSS.t57 208.07
R132 VSS.n74 VSS.n73 199.794
R133 VSS.n77 VSS.n12 199.794
R134 VSS VSS.n10 199.794
R135 VSS VSS.n8 199.794
R136 VSS VSS.n1 199.794
R137 VSS.n28 VSS.n27 199.794
R138 VSS.n32 VSS.n31 199.794
R139 VSS.n63 VSS.n50 164.93
R140 VSS.n47 VSS.n19 164.93
R141 VSS.n68 VSS.n16 164.93
R142 VSS.n57 VSS.n16 164.93
R143 VSS.n39 VSS.n18 164.93
R144 VSS.n25 VSS.n18 164.93
R145 VSS.n40 VSS.t12 106.218
R146 VSS.n24 VSS.t55 106.218
R147 VSS.n67 VSS.t57 104.763
R148 VSS.n64 VSS.t56 104.763
R149 VSS.n58 VSS.t56 104.763
R150 VSS.n48 VSS.t12 103.308
R151 VSS.n73 VSS.t9 82.8576
R152 VSS.n12 VSS.t17 82.8576
R153 VSS.n10 VSS.t15 82.8576
R154 VSS.n8 VSS.t36 82.8576
R155 VSS.n1 VSS.t24 82.8576
R156 VSS.n27 VSS.t21 82.8576
R157 VSS.n31 VSS.t47 82.8576
R158 VSS.n73 VSS.t38 81.4291
R159 VSS.n12 VSS.t30 81.4291
R160 VSS.n10 VSS.t28 81.4291
R161 VSS.n8 VSS.t34 81.4291
R162 VSS.n1 VSS.t22 81.4291
R163 VSS.n27 VSS.t19 81.4291
R164 VSS.n31 VSS.t43 81.4291
R165 VSS.n66 VSS.t0 65.4767
R166 VSS.n49 VSS.n48 64.0217
R167 VSS.t50 VSS.n17 64.0217
R168 VSS.n65 VSS.n64 64.0217
R169 VSS.n41 VSS.n19 62.4724
R170 VSS.n59 VSS.n50 62.4724
R171 VSS.n49 VSS.t50 40.7412
R172 VSS.n24 VSS.n17 40.7412
R173 VSS.n67 VSS.n66 40.7412
R174 VSS.t0 VSS.n65 39.2862
R175 VSS.n62 VSS.n61 10.7168
R176 VSS.n61 VSS.n60 10.7168
R177 VSS.n42 VSS.n20 10.7168
R178 VSS.n46 VSS.n20 10.7168
R179 VSS.n69 VSS.n15 10.7168
R180 VSS.n56 VSS.n15 10.7168
R181 VSS.n38 VSS.n23 10.7168
R182 VSS.n26 VSS.n23 10.7168
R183 VSS.n62 VSS.n51 9.3005
R184 VSS.n61 VSS.n52 9.3005
R185 VSS.n60 VSS.n53 9.3005
R186 VSS.n44 VSS.n20 9.3005
R187 VSS.n46 VSS.n45 9.3005
R188 VSS.n43 VSS.n42 9.3005
R189 VSS.n15 VSS.n14 9.3005
R190 VSS.n56 VSS.n55 9.3005
R191 VSS.n70 VSS.n69 9.3005
R192 VSS.n36 VSS.n23 9.3005
R193 VSS.n35 VSS.n26 9.3005
R194 VSS.n38 VSS.n37 9.3005
R195 VSS.n54 VSS.n53 5.56717
R196 VSS.n43 VSS.n22 5.56717
R197 VSS.n37 VSS.n22 5.41717
R198 VSS.n51 VSS.n13 5.41717
R199 VSS.n45 VSS.n21 5.41717
R200 VSS.n71 VSS.n70 5.41717
R201 VSS.n55 VSS.n54 5.41717
R202 VSS.n35 VSS.n34 5.41717
R203 VSS.n78 VSS.n77 3.43911
R204 VSS.n28 VSS.n5 3.43911
R205 VSS.n3 VSS.n0 3.4105
R206 VSS VSS.n85 3.4105
R207 VSS.n4 VSS.n2 3.4105
R208 VSS VSS.n6 3.4105
R209 VSS.n81 VSS.n9 3.4105
R210 VSS.n80 VSS 3.4105
R211 VSS.n79 VSS.n11 3.4105
R212 VSS.n85 VSS.n84 3.4105
R213 VSS.n83 VSS.n4 3.4105
R214 VSS VSS.n6 3.4105
R215 VSS.n82 VSS.n81 3.4105
R216 VSS.n80 VSS.n7 3.4105
R217 VSS.t48 VSS.t1 2.91055
R218 VSS.n84 VSS.n5 1.73427
R219 VSS.n78 VSS.n7 1.73427
R220 VSS.t45 VSS.t13 1.45553
R221 VSS.t42 VSS.t58 1.45553
R222 VSS.t44 VSS.t46 1.45553
R223 VSS.t4 VSS.t25 1.45553
R224 VSS.t2 VSS.t10 1.45553
R225 VSS.t39 VSS.t23 1.45553
R226 VSS.t31 VSS.t52 1.45553
R227 VSS.t37 VSS.t41 1.45553
R228 VSS.t51 VSS.t8 1.45553
R229 VSS.t6 VSS.t3 1.45553
R230 VSS.n33 VSS.n32 0.3005
R231 VSS.n74 VSS.n72 0.3005
R232 VSS.n22 VSS.n21 0.1505
R233 VSS.n34 VSS.n21 0.1505
R234 VSS.n34 VSS.n33 0.1505
R235 VSS.n32 VSS.n30 0.1505
R236 VSS.n30 VSS.n29 0.1505
R237 VSS.n29 VSS.n28 0.1505
R238 VSS.n28 VSS.n0 0.1505
R239 VSS VSS.n0 0.1505
R240 VSS VSS.n2 0.1505
R241 VSS VSS.n2 0.1505
R242 VSS.n9 VSS 0.1505
R243 VSS VSS.n9 0.1505
R244 VSS.n11 VSS 0.1505
R245 VSS.n77 VSS.n11 0.1505
R246 VSS.n77 VSS.n76 0.1505
R247 VSS.n76 VSS.n75 0.1505
R248 VSS.n75 VSS.n74 0.1505
R249 VSS.n72 VSS.n71 0.1505
R250 VSS.n71 VSS.n13 0.1505
R251 VSS.n54 VSS.n13 0.1505
R252 VSS.n52 VSS.n51 0.105151
R253 VSS.n53 VSS.n52 0.105151
R254 VSS.n44 VSS.n43 0.105151
R255 VSS.n45 VSS.n44 0.105151
R256 VSS.n70 VSS.n14 0.105151
R257 VSS.n55 VSS.n14 0.105151
R258 VSS.n37 VSS.n36 0.105151
R259 VSS.n36 VSS.n35 0.105151
R260 VSS.n85 VSS.n3 0.0569
R261 VSS.n85 VSS.n4 0.0569
R262 VSS.n6 VSS.n4 0.0569
R263 VSS.n81 VSS.n6 0.0569
R264 VSS.n81 VSS.n80 0.0569
R265 VSS.n80 VSS.n79 0.0569
R266 VSS.n84 VSS.n83 0.03434
R267 VSS.n83 VSS 0.03434
R268 VSS VSS.n82 0.03434
R269 VSS.n82 VSS.n7 0.03434
R270 VSS.n5 VSS.n3 0.0288317
R271 VSS.n79 VSS.n78 0.0288317
R272 Di_n Di_n.n2 603.328
R273 Di_n.n1 Di_n.t14 164.137
R274 Di_n.n1 Di_n.t12 164.137
R275 Di_n.n0 Di_n.t13 164.137
R276 Di_n.n0 Di_n.t15 164.137
R277 Di_n.n2 Di_n.t4 133.679
R278 Di_n.n2 Di_n.t3 131.333
R279 Di_n.n11 Di_n.n9 102.382
R280 Di_n.n4 Di_n.n3 101.79
R281 Di_n.n6 Di_n.n5 101.79
R282 Di_n.n8 Di_n.n7 101.79
R283 Di_n.n11 Di_n.n10 101.79
R284 Di_n Di_n.n0 73.6595
R285 Di_n.n13 Di_n.n1 73.3637
R286 Di_n.n3 Di_n.t6 40.7148
R287 Di_n.n5 Di_n.t11 40.7148
R288 Di_n.n7 Di_n.t8 40.7148
R289 Di_n.n10 Di_n.t10 40.7148
R290 Di_n.n9 Di_n.t9 40.7148
R291 Di_n.n3 Di_n.t1 40.0005
R292 Di_n.n5 Di_n.t7 40.0005
R293 Di_n.n7 Di_n.t5 40.0005
R294 Di_n.n10 Di_n.t2 40.0005
R295 Di_n.n9 Di_n.t0 40.0005
R296 Di_n.n13 Di_n.n12 8.49997
R297 Di_n.n4 Di_n 4.4346
R298 Di_n.n8 Di_n.n6 0.592167
R299 Di_n.n6 Di_n.n4 0.592167
R300 Di_n Di_n.n13 0.283833
R301 Di_n.n12 Di_n.n11 0.279667
R302 Di_n.n12 Di_n.n8 0.279667
R303 Vout_p Vout_p.n2 602.75
R304 Vout_p.n6 Vout_p.n4 199.486
R305 Vout_p.n7 Vout_p.n3 198.894
R306 Vout_p.n6 Vout_p.n5 198.894
R307 Vout_p.n0 Vout_p.t9 164.137
R308 Vout_p.n0 Vout_p.t10 164.137
R309 Vout_p.n1 Vout_p.t11 164.137
R310 Vout_p.n1 Vout_p.t8 164.137
R311 Vout_p.n2 Vout_p.t4 133.679
R312 Vout_p.n2 Vout_p.t5 131.333
R313 Vout_p.n3 Vout_p.t7 81.4291
R314 Vout_p.n5 Vout_p.t2 81.4291
R315 Vout_p.n4 Vout_p.t3 81.4291
R316 Vout_p.n3 Vout_p.t6 80.0005
R317 Vout_p.n5 Vout_p.t0 80.0005
R318 Vout_p.n4 Vout_p.t1 80.0005
R319 Vout_p Vout_p.n0 77.2722
R320 Vout_p.n9 Vout_p.n1 77.1531
R321 Vout_p Vout_p.n8 3.84383
R322 Vout_p.n9 Vout_p 3.84383
R323 Vout_p.n8 Vout_p.n7 3.73637
R324 Vout_p.n7 Vout_p.n6 1.17967
R325 Vout_p.n8 Vout_p 0.107033
R326 Vout_p Vout_p.n9 0.107033
R327 Vin_p.n3 Vin_p.t6 231.618
R328 Vin_p.n5 Vin_p.t9 231.618
R329 Vin_p.n4 Vin_p.t2 231.618
R330 Vin_p.n1 Vin_p.t8 231.618
R331 Vin_p.n0 Vin_p.t3 231.618
R332 Vin_p.n3 Vin_p.t7 231.618
R333 Vin_p.n5 Vin_p.t0 231.618
R334 Vin_p.n4 Vin_p.t4 231.618
R335 Vin_p.n1 Vin_p.t1 231.618
R336 Vin_p.n0 Vin_p.t5 231.618
R337 Vin_p.n6 Vin_p.n4 73.9026
R338 Vin_p.n2 Vin_p.n0 73.9026
R339 Vin_p Vin_p.n3 73.311
R340 Vin_p.n6 Vin_p.n5 73.311
R341 Vin_p.n2 Vin_p.n1 73.311
R342 Vin_p Vin_p.n6 0.592167
R343 Vin_p Vin_p.n2 0.592167
R344 Vin_n.n3 Vin_n.t1 231.618
R345 Vin_n.n5 Vin_n.t7 231.618
R346 Vin_n.n4 Vin_n.t2 231.618
R347 Vin_n.n1 Vin_n.t6 231.618
R348 Vin_n.n0 Vin_n.t3 231.618
R349 Vin_n.n3 Vin_n.t4 231.618
R350 Vin_n.n5 Vin_n.t8 231.618
R351 Vin_n.n4 Vin_n.t0 231.618
R352 Vin_n.n1 Vin_n.t9 231.618
R353 Vin_n.n0 Vin_n.t5 231.618
R354 Vin_n.n6 Vin_n.n4 73.9026
R355 Vin_n.n2 Vin_n.n0 73.9026
R356 Vin_n Vin_n.n3 73.311
R357 Vin_n.n6 Vin_n.n5 73.311
R358 Vin_n.n2 Vin_n.n1 73.311
R359 Vin_n Vin_n.n6 0.592167
R360 Vin_n Vin_n.n2 0.592167
R361 Di_p Di_p.n4 603.328
R362 Di_p.n0 Di_p.t14 164.137
R363 Di_p.n0 Di_p.t12 164.137
R364 Di_p.n13 Di_p.t15 164.137
R365 Di_p.n13 Di_p.t13 164.137
R366 Di_p.n4 Di_p.t1 133.679
R367 Di_p.n4 Di_p.t0 131.333
R368 Di_p.n3 Di_p.n1 102.382
R369 Di_p.n6 Di_p.n5 101.79
R370 Di_p.n8 Di_p.n7 101.79
R371 Di_p.n10 Di_p.n9 101.79
R372 Di_p.n3 Di_p.n2 101.79
R373 Di_p Di_p.n13 73.6595
R374 Di_p.n12 Di_p.n0 73.3637
R375 Di_p.n5 Di_p.t9 40.7148
R376 Di_p.n7 Di_p.t4 40.7148
R377 Di_p.n9 Di_p.t10 40.7148
R378 Di_p.n2 Di_p.t5 40.7148
R379 Di_p.n1 Di_p.t8 40.7148
R380 Di_p.n5 Di_p.t11 40.0005
R381 Di_p.n7 Di_p.t3 40.0005
R382 Di_p.n9 Di_p.t7 40.0005
R383 Di_p.n2 Di_p.t2 40.0005
R384 Di_p.n1 Di_p.t6 40.0005
R385 Di_p.n12 Di_p.n11 8.49997
R386 Di_p.n6 Di_p 4.4346
R387 Di_p.n10 Di_p.n8 0.592167
R388 Di_p.n8 Di_p.n6 0.592167
R389 Di_p Di_p.n12 0.283833
R390 Di_p.n11 Di_p.n3 0.279667
R391 Di_p.n11 Di_p.n10 0.279667
R392 Vout_n.n4 Vout_n.n0 602.63
R393 Vout_n.n7 Vout_n.n5 199.486
R394 Vout_n.n9 Vout_n.n8 198.894
R395 Vout_n.n7 Vout_n.n6 198.894
R396 Vout_n.n1 Vout_n.t10 164.137
R397 Vout_n.n1 Vout_n.t11 164.137
R398 Vout_n.n2 Vout_n.t8 164.137
R399 Vout_n.n2 Vout_n.t9 164.137
R400 Vout_n.n0 Vout_n.t0 133.679
R401 Vout_n.n0 Vout_n.t1 131.333
R402 Vout_n.n8 Vout_n.t2 81.4291
R403 Vout_n.n6 Vout_n.t6 81.4291
R404 Vout_n.n5 Vout_n.t5 81.4291
R405 Vout_n.n8 Vout_n.t3 80.0005
R406 Vout_n.n6 Vout_n.t4 80.0005
R407 Vout_n.n5 Vout_n.t7 80.0005
R408 Vout_n Vout_n.n2 77.2722
R409 Vout_n.n3 Vout_n.n1 77.1531
R410 Vout_n Vout_n.n9 3.85543
R411 Vout_n Vout_n.n3 3.84383
R412 Vout_n.n4 Vout_n 3.84383
R413 Vout_n.n9 Vout_n.n7 1.17967
R414 Vout_n.n3 Vout_n 0.107033
R415 Vout_n Vout_n.n4 0.107033
R416 CLK_bar.n8 CLK_bar.t5 231.618
R417 CLK_bar.n6 CLK_bar.t4 231.618
R418 CLK_bar.n5 CLK_bar.t2 231.618
R419 CLK_bar.n3 CLK_bar.t3 231.618
R420 CLK_bar.n1 CLK_bar.t8 231.618
R421 CLK_bar.n0 CLK_bar.t10 231.618
R422 CLK_bar.n8 CLK_bar.t1 231.618
R423 CLK_bar.n6 CLK_bar.t0 231.618
R424 CLK_bar.n5 CLK_bar.t11 231.618
R425 CLK_bar.n3 CLK_bar.t7 231.618
R426 CLK_bar.n1 CLK_bar.t9 231.618
R427 CLK_bar.n0 CLK_bar.t6 231.618
R428 CLK_bar.n7 CLK_bar.n5 73.9026
R429 CLK_bar.n2 CLK_bar.n0 73.9026
R430 CLK_bar.n9 CLK_bar.n8 73.311
R431 CLK_bar.n7 CLK_bar.n6 73.311
R432 CLK_bar.n4 CLK_bar.n3 73.311
R433 CLK_bar.n2 CLK_bar.n1 73.311
R434 CLK_bar.n9 CLK_bar.n7 0.592167
R435 CLK_bar.n4 CLK_bar.n2 0.592167
R436 CLK_bar CLK_bar.n9 0.296333
R437 CLK_bar CLK_bar.n4 0.296333
R438 VDD.n18 VDD.t5 735.818
R439 VDD.n59 VDD.t11 735.818
R440 VDD.n20 VDD.t7 733.472
R441 VDD.n53 VDD.t9 733.472
R442 VDD.n81 VDD.t23 370.702
R443 VDD.n105 VDD.t30 369.529
R444 VDD.n66 VDD.t22 340.228
R445 VDD.n116 VDD.t29 339.286
R446 VDD.n103 VDD.n34 302.69
R447 VDD.n97 VDD.n96 302.69
R448 VDD VDD.n39 302.69
R449 VDD.n90 VDD.n89 302.69
R450 VDD.n87 VDD.n44 302.69
R451 VDD.n9 VDD.t4 204.514
R452 VDD.n7 VDD.t8 203.571
R453 VDD.n117 VDD.n116 187.567
R454 VDD.n66 VDD.n64 187.567
R455 VDD.n118 VDD.n117 140.934
R456 VDD.n70 VDD.n64 140.934
R457 VDD.n8 VDD.n7 135.714
R458 VDD.n9 VDD.n8 135.714
R459 VDD.t12 VDD.t29 134.773
R460 VDD.t22 VDD.t14 134.773
R461 VDD.t8 VDD.t10 134.773
R462 VDD.t4 VDD.t6 134.773
R463 VDD.t25 VDD.t12 102.728
R464 VDD.t14 VDD.t16 102.257
R465 VDD.n115 VDD.n114 92.5005
R466 VDD.n116 VDD.n115 92.5005
R467 VDD.n27 VDD.n26 92.5005
R468 VDD.n68 VDD.n67 92.5005
R469 VDD.n67 VDD.n66 92.5005
R470 VDD.n69 VDD.n65 92.5005
R471 VDD.n11 VDD.n10 92.5005
R472 VDD.n10 VDD.n9 92.5005
R473 VDD.n3 VDD.n2 92.5005
R474 VDD.n8 VDD.n3 92.5005
R475 VDD.n6 VDD.n5 92.5005
R476 VDD.n7 VDD.n6 92.5005
R477 VDD.n115 VDD.n27 86.4005
R478 VDD.n67 VDD.n65 86.4005
R479 VDD.n6 VDD.n3 86.4005
R480 VDD.n10 VDD.n3 86.4005
R481 VDD.t27 VDD.t31 68.3289
R482 VDD.n34 VDD.t13 68.0124
R483 VDD.n96 VDD.t34 68.0124
R484 VDD.n39 VDD.t32 68.0124
R485 VDD.n89 VDD.t21 68.0124
R486 VDD.n44 VDD.t17 68.0124
R487 VDD.t16 VDD.t18 67.3864
R488 VDD.t1 VDD.t0 67.3864
R489 VDD.t20 VDD.t27 67.3864
R490 VDD.t31 VDD.t3 67.3864
R491 VDD.t3 VDD.t2 67.3864
R492 VDD.t33 VDD.t25 67.3864
R493 VDD.n34 VDD.t26 66.8398
R494 VDD.n96 VDD.t24 66.8398
R495 VDD.n39 VDD.t28 66.8398
R496 VDD.n89 VDD.t19 66.8398
R497 VDD.n44 VDD.t15 66.8398
R498 VDD.n117 VDD.n27 19.6319
R499 VDD.n65 VDD.n64 19.6319
R500 VDD.n114 VDD.n26 9.2165
R501 VDD.n118 VDD.n26 9.2165
R502 VDD.n70 VDD.n69 9.2165
R503 VDD.n69 VDD.n68 9.2165
R504 VDD.n5 VDD.n2 9.2165
R505 VDD.n11 VDD.n2 9.2165
R506 VDD.n72 VDD.n71 5.12967
R507 VDD.n120 VDD.n119 5.12967
R508 VDD.n113 VDD.n112 5.12967
R509 VDD.n79 VDD.n49 5.12967
R510 VDD.n4 VDD.n0 5.12967
R511 VDD.n13 VDD.n12 5.12967
R512 VDD.n114 VDD.n113 4.6505
R513 VDD.n26 VDD.n25 4.6505
R514 VDD.n119 VDD.n118 4.6505
R515 VDD.n69 VDD.n63 4.6505
R516 VDD.n68 VDD.n49 4.6505
R517 VDD.n71 VDD.n70 4.6505
R518 VDD.n2 VDD.n1 4.6505
R519 VDD.n12 VDD.n11 4.6505
R520 VDD.n5 VDD.n4 4.6505
R521 VDD.n73 VDD.n62 3.43958
R522 VDD.n122 VDD.n121 3.43958
R523 VDD.n61 VDD.n60 3.43958
R524 VDD.n123 VDD.n21 3.43958
R525 VDD.n30 VDD.n24 3.4105
R526 VDD.n50 VDD.n48 3.4105
R527 VDD.n79 VDD.n78 3.4105
R528 VDD.n80 VDD.n47 3.4105
R529 VDD.n82 VDD.n81 3.4105
R530 VDD.n45 VDD.n43 3.4105
R531 VDD.n87 VDD.n86 3.4105
R532 VDD.n88 VDD.n42 3.4105
R533 VDD.n91 VDD.n90 3.4105
R534 VDD.n40 VDD.n38 3.4105
R535 VDD VDD.n94 3.4105
R536 VDD.n95 VDD.n37 3.4105
R537 VDD.n98 VDD.n97 3.4105
R538 VDD.n35 VDD.n33 3.4105
R539 VDD.n103 VDD.n102 3.4105
R540 VDD.n104 VDD.n32 3.4105
R541 VDD.n106 VDD.n105 3.4105
R542 VDD.n29 VDD.n28 3.4105
R543 VDD.n112 VDD.n111 3.4105
R544 VDD.n58 VDD.n57 3.4105
R545 VDD.n54 VDD.n53 3.4105
R546 VDD.n14 VDD.n0 3.4105
R547 VDD VDD.n131 3.4105
R548 VDD.n15 VDD.n13 3.4105
R549 VDD.n127 VDD.n18 3.4105
R550 VDD.n126 VDD.n19 3.4105
R551 VDD.n52 VDD.n51 3.4105
R552 VDD.n57 VDD.n56 3.4105
R553 VDD.n55 VDD.n54 3.4105
R554 VDD.n16 VDD.n14 3.4105
R555 VDD.n131 VDD.n130 3.4105
R556 VDD.n129 VDD.n15 3.4105
R557 VDD.n128 VDD.n127 3.4105
R558 VDD.n126 VDD.n17 3.4105
R559 VDD.n125 VDD.n124 3.4105
R560 VDD.n109 VDD.n30 3.4105
R561 VDD.n23 VDD.n22 3.4105
R562 VDD.n75 VDD.n74 3.4105
R563 VDD.n76 VDD.n50 3.4105
R564 VDD.n78 VDD.n77 3.4105
R565 VDD.n47 VDD.n46 3.4105
R566 VDD.n83 VDD.n82 3.4105
R567 VDD.n84 VDD.n45 3.4105
R568 VDD.n86 VDD.n85 3.4105
R569 VDD.n42 VDD.n41 3.4105
R570 VDD.n92 VDD.n91 3.4105
R571 VDD.n93 VDD.n40 3.4105
R572 VDD.n94 VDD 3.4105
R573 VDD.n37 VDD.n36 3.4105
R574 VDD.n99 VDD.n98 3.4105
R575 VDD.n100 VDD.n35 3.4105
R576 VDD.n102 VDD.n101 3.4105
R577 VDD.n32 VDD.n31 3.4105
R578 VDD.n107 VDD.n106 3.4105
R579 VDD.n108 VDD.n29 3.4105
R580 VDD.n111 VDD.n110 3.4105
R581 VDD.n123 VDD.n122 1.76571
R582 VDD.n62 VDD.n61 1.76571
R583 VDD.n73 VDD.n72 1.72871
R584 VDD.n121 VDD.n120 1.72871
R585 VDD.n60 VDD.n59 1.72871
R586 VDD.n21 VDD.n20 1.72871
R587 VDD.t2 VDD.t33 0.94296
R588 VDD.t18 VDD.t1 0.47173
R589 VDD.t0 VDD.t20 0.47173
R590 VDD.n72 VDD.n48 0.1505
R591 VDD.n79 VDD.n48 0.1505
R592 VDD.n80 VDD.n79 0.1505
R593 VDD.n81 VDD.n80 0.1505
R594 VDD.n81 VDD.n43 0.1505
R595 VDD.n87 VDD.n43 0.1505
R596 VDD.n88 VDD.n87 0.1505
R597 VDD.n90 VDD.n88 0.1505
R598 VDD.n90 VDD.n38 0.1505
R599 VDD VDD.n38 0.1505
R600 VDD.n95 VDD 0.1505
R601 VDD.n97 VDD.n95 0.1505
R602 VDD.n97 VDD.n33 0.1505
R603 VDD.n103 VDD.n33 0.1505
R604 VDD.n104 VDD.n103 0.1505
R605 VDD.n105 VDD.n104 0.1505
R606 VDD.n105 VDD.n28 0.1505
R607 VDD.n112 VDD.n28 0.1505
R608 VDD.n112 VDD.n24 0.1505
R609 VDD.n120 VDD.n24 0.1505
R610 VDD.n59 VDD.n58 0.1505
R611 VDD.n58 VDD.n53 0.1505
R612 VDD.n53 VDD.n0 0.1505
R613 VDD VDD.n0 0.1505
R614 VDD VDD.n13 0.1505
R615 VDD.n18 VDD.n13 0.1505
R616 VDD.n19 VDD.n18 0.1505
R617 VDD.n20 VDD.n19 0.1505
R618 VDD.n113 VDD.n25 0.0905
R619 VDD.n119 VDD.n25 0.0905
R620 VDD.n71 VDD.n63 0.0905
R621 VDD.n63 VDD.n49 0.0905
R622 VDD.n4 VDD.n1 0.0905
R623 VDD.n12 VDD.n1 0.0905
R624 VDD.n74 VDD.n50 0.0569
R625 VDD.n78 VDD.n50 0.0569
R626 VDD.n78 VDD.n47 0.0569
R627 VDD.n82 VDD.n47 0.0569
R628 VDD.n82 VDD.n45 0.0569
R629 VDD.n86 VDD.n45 0.0569
R630 VDD.n86 VDD.n42 0.0569
R631 VDD.n91 VDD.n42 0.0569
R632 VDD.n91 VDD.n40 0.0569
R633 VDD.n94 VDD.n40 0.0569
R634 VDD.n94 VDD.n37 0.0569
R635 VDD.n98 VDD.n37 0.0569
R636 VDD.n98 VDD.n35 0.0569
R637 VDD.n102 VDD.n35 0.0569
R638 VDD.n102 VDD.n32 0.0569
R639 VDD.n106 VDD.n32 0.0569
R640 VDD.n106 VDD.n29 0.0569
R641 VDD.n111 VDD.n29 0.0569
R642 VDD.n111 VDD.n30 0.0569
R643 VDD.n30 VDD.n23 0.0569
R644 VDD.n57 VDD.n52 0.0569
R645 VDD.n57 VDD.n54 0.0569
R646 VDD.n54 VDD.n14 0.0569
R647 VDD.n131 VDD.n14 0.0569
R648 VDD.n131 VDD.n15 0.0569
R649 VDD.n127 VDD.n15 0.0569
R650 VDD.n127 VDD.n126 0.0569
R651 VDD.n126 VDD.n125 0.0569
R652 VDD.n61 VDD.n51 0.03434
R653 VDD.n56 VDD.n51 0.03434
R654 VDD.n56 VDD.n55 0.03434
R655 VDD.n55 VDD.n16 0.03434
R656 VDD.n130 VDD.n16 0.03434
R657 VDD.n130 VDD.n129 0.03434
R658 VDD.n129 VDD.n128 0.03434
R659 VDD.n128 VDD.n17 0.03434
R660 VDD.n124 VDD.n17 0.03434
R661 VDD.n124 VDD.n123 0.03434
R662 VDD.n75 VDD.n62 0.03434
R663 VDD.n76 VDD.n75 0.03434
R664 VDD.n77 VDD.n76 0.03434
R665 VDD.n77 VDD.n46 0.03434
R666 VDD.n83 VDD.n46 0.03434
R667 VDD.n84 VDD.n83 0.03434
R668 VDD.n85 VDD.n84 0.03434
R669 VDD.n85 VDD.n41 0.03434
R670 VDD.n92 VDD.n41 0.03434
R671 VDD.n93 VDD.n92 0.03434
R672 VDD VDD.n93 0.03434
R673 VDD VDD.n36 0.03434
R674 VDD.n99 VDD.n36 0.03434
R675 VDD.n100 VDD.n99 0.03434
R676 VDD.n101 VDD.n100 0.03434
R677 VDD.n101 VDD.n31 0.03434
R678 VDD.n107 VDD.n31 0.03434
R679 VDD.n108 VDD.n107 0.03434
R680 VDD.n110 VDD.n108 0.03434
R681 VDD.n110 VDD.n109 0.03434
R682 VDD.n109 VDD.n22 0.03434
R683 VDD.n122 VDD.n22 0.03434
R684 VDD.n121 VDD.n23 0.0283716
R685 VDD.n74 VDD.n73 0.0283716
R686 VDD.n60 VDD.n52 0.0283716
R687 VDD.n125 VDD.n21 0.0283716
C0 VDD latch.inv0.VDD 3.97f
.ends






































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































* expanding   symbol:  RS_latch.sym # of pins=5
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/RS_latch.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/RS_latch.sch
.subckt RS_latch VDD R Q S Q_bar
*.iopin VDD
*.opin Q
*.opin Q_bar
*.ipin R
*.ipin S
x1 VDD R Q_bar Q nor
x2 VDD Q S Q_bar nor
.ends


* expanding   symbol:  nor.sym # of pins=4
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/nor.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/nor.sch
.subckt nor VDD A B out
*.iopin VDD
*.ipin A
*.ipin B
*.opin out
XM1 out B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out B net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
**** begin user architecture code

.model filesrc filesource (file="staircase_voltage.txt" amploffset=[Vcm] amplscale=[1] timeoffset=0
+ timescale=1 timerelative=false amplstep=false)

**** end user architecture code
.end

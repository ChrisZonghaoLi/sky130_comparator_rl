* transient analysis clk-2-Q
*tran 1p 3n
*plot v(Vclk) v(Vclk_bar)
*plot v(Vout_n) v(Vout_p)
*plot v(Di_p) v(Di_n)
*plot v(Q) v(Q_bar)
*wrdata double_tail_comp_tb_Voutn Vout_n 
*wrdata double_tail_comp_tb_Voutp Vout_p 
*wrdata double_tail_comp_tb_Vclk Vclk

* power consumption
*plot @Rdummy[i]
*wrdata double_tail_comp_tb_Ibias @Rdummy[i]

* kickback noise
*plot {Vp_kn-Vn_kn}
*wrdata double_tail_comp_tb_Vn_kn Vn_kn 
*wrdata double_tail_comp_tb_Vp_kn Vp_kn 

* metastability
*plot {Vout_p_ms-Vout_n_ms}
*wrdata double_tail_comp_tb_Voutn_ms Vout_n_ms 
*wrdata double_tail_comp_tb_Voutp_ms Vout_p_ms 

* op analysis
alter Vclk dc=1.8
alter Vclk_bar dc=0
alter Vdiff dc=0
op
.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/comparator_transfer_learning/pex/simulations/double_tail_comp_tb_dev_params.spice

magic
tech sky130A
magscale 1 2
timestamp 1706304417
<< pwell >>
rect -92 443 236 599
<< nmos >>
rect 57 479 87 563
<< ndiff >>
rect -56 541 57 563
rect -56 501 -20 541
rect 20 501 57 541
rect -56 479 57 501
rect 87 541 200 563
rect 87 501 124 541
rect 164 501 200 541
rect 87 479 200 501
<< ndiffc >>
rect -20 501 20 541
rect 124 501 164 541
<< poly >>
rect 32 659 112 679
rect 32 619 52 659
rect 92 619 112 659
rect 32 599 112 619
rect 57 563 87 599
rect 57 443 87 479
<< polycont >>
rect 52 619 92 659
<< locali >>
rect 32 659 112 679
rect 32 619 52 659
rect 92 619 112 659
rect 32 599 112 619
rect -30 541 30 557
rect -30 501 -20 541
rect 20 501 30 541
rect -30 485 30 501
rect 114 541 174 557
rect 114 501 124 541
rect 164 501 174 541
rect 114 485 174 501
<< viali >>
rect 52 619 92 659
rect -20 501 20 541
rect 124 501 164 541
<< metal1 >>
rect 32 659 112 679
rect 32 619 52 659
rect 92 619 112 659
rect 32 599 112 619
rect -30 541 30 557
rect -30 501 -20 541
rect 20 501 30 541
rect -30 329 30 501
rect 114 541 174 557
rect 114 501 124 541
rect 164 501 174 541
rect 114 329 174 501
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1706648821
<< nwell >>
rect -92 132 380 684
<< pmos >>
rect 57 437 87 521
rect 200 437 230 521
<< pdiff >>
rect -56 499 57 521
rect -56 459 -20 499
rect 20 459 57 499
rect -56 437 57 459
rect 87 499 200 521
rect 87 459 124 499
rect 164 459 200 499
rect 87 437 200 459
rect 230 499 343 521
rect 230 459 268 499
rect 308 459 343 499
rect 230 437 343 459
<< pdiffc >>
rect -20 459 20 499
rect 124 459 164 499
rect 268 459 308 499
<< poly >>
rect 57 617 230 637
rect 57 577 77 617
rect 117 577 170 617
rect 210 577 230 617
rect 57 557 230 577
rect 57 521 87 557
rect 200 521 230 557
rect 57 401 87 437
rect 200 401 230 437
<< polycont >>
rect 77 577 117 617
rect 170 577 210 617
<< locali >>
rect 57 617 230 637
rect 57 577 77 617
rect 117 577 170 617
rect 210 577 230 617
rect 57 557 230 577
rect -30 499 30 515
rect -30 459 -20 499
rect 20 459 30 499
rect -30 443 30 459
rect 114 499 174 515
rect 114 459 124 499
rect 164 459 174 499
rect 114 443 174 459
rect 258 499 318 515
rect 258 459 268 499
rect 308 459 318 499
rect 258 443 318 459
<< viali >>
rect 77 577 117 617
rect 170 577 210 617
rect -20 459 20 499
rect 124 459 164 499
rect 268 459 308 499
<< metal1 >>
rect 57 617 230 757
rect 57 577 77 617
rect 117 577 170 617
rect 210 577 230 617
rect 57 557 230 577
rect -30 499 30 515
rect -30 459 -20 499
rect 20 459 30 499
rect -30 227 30 459
rect 114 499 174 515
rect 114 459 124 499
rect 164 459 174 499
rect 114 227 174 459
rect 258 499 318 515
rect 258 459 268 499
rect 308 459 318 499
rect 258 227 318 459
<< end >>

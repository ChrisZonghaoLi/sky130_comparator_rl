magic
tech sky130A
timestamp 1709070663
<< via4 >>
rect -60 -60 60 60
<< metal5 >>
rect -100 60 100 100
rect -100 -60 -60 60
rect 60 -60 100 60
rect -100 -100 100 -60
<< end >>

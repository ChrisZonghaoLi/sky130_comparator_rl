** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp_pex_tb.sch
**.subckt double_tail_comp_pex_tb Di_n Di_p Vout_n Vout_p Q Q_bar Di_n_mc Di_p_mc Vout_n_mc
*+ Vout_p_mc Di_n_ms Di_p_ms Vout_n_ms Vout_p_ms Di_n_kn Di_p_kn Vout_n_kn Vout_p_kn
*.opin Di_n
*.opin Di_p
*.opin Vout_n
*.opin Vout_p
*.opin Q
*.opin Q_bar
*.opin Di_n_mc
*.opin Di_p_mc
*.opin Vout_n_mc
*.opin Vout_p_mc
*.opin Di_n_ms
*.opin Di_p_ms
*.opin Vout_n_ms
*.opin Vout_p_ms
*.opin Di_n_kn
*.opin Di_p_kn
*.opin Vout_n_kn
*.opin Vout_p_kn
x1 net1 Vclk_bar Vout_n Vout_p Di_n Di_p Vcm net10 Vclk GND double_tail_comp
VDD net1 net9 VDD
Vclk Vclk GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar Vclk_bar GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm Vcm GND dc Vcm
Vdiff net10 Vcm dc Vin
C2 Q_bar GND 10f m=1
C3 Q GND 10f m=1
x2 net17 Vout_n Q Vout_p Q_bar RS_latch
x3 net4 net3 Vout_n_mc Vout_p_mc Di_n_mc Di_p_mc net2 Vsc net15 GND double_tail_comp
VDD2 net4 GND VDD
Vclk2 net15 GND PULSE(0 VDD 0 Tr Tf Tclk_pk Tclk 0)
Vclk_bar2 net3 GND PULSE(0 VDD Tclk_pk Tr Tf Tclk_pk Tclk 0)
Vcm2 net2 GND dc Vcm
ASRC1 %v([ Vsc ]) filesrc
x4 net8 net7 Vout_n_ms Vout_p_ms Di_n_ms Di_p_ms net5 net6 net16 GND double_tail_comp
VDD3 net8 GND VDD
Vclk3 net16 GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar3 net7 GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm3 net5 GND dc Vcm
Vdiff2 net6 net5 dc Vin_min
VDD_latch net17 GND VDD
Rdummy net9 GND 1 m=1
x5 net13 net12 Vout_n_kn Vout_p_kn Di_n_kn Di_p_kn Vn_kn Vp_kn net18 GND double_tail_comp
VDD4 net13 GND VDD
Vclk4 net18 GND PULSE(0 VDD Tdelay Tr Tf Tclk_pk Tclk 0)
Vclk_bar5 net12 GND PULSE(0 VDD Tdelay_bar Tr Tf Tclk_pk Tclk 0)
Vcm4 net11 GND dc Vcm
Vdiff4 net14 net11 dc Vin
Rdummyn net11 Vn_kn 8k m=1
Rdummyp net14 Vp_kn 8k m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /usr/local/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



*.OPTIONS maxord=1
*.OPTIONS itl1=200
*.OPTIONS itl2=200
*.OPTIONS itl4=200

* save all voltage and current
.save all
.options savecurrents
.options seed=random

.control
set filetype=ascii
set units=degrees

* RC extracted comparator netlist
.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/sky130_comparator/netgen/double_tail/TCL/double_tail_comparator_pex.spice
* analyses
.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/sky130_comparator/xschem/simulations/double_tail_comp_pex_tb_analyses.spice
* stimulus variables
.include /autofs/fs1.ece/fs1.eecg.tcc/lizongh2/sky130_comparator/xschem/simulations/double_tail_comp_pex_tb_vars.spice

.endc


**** end user architecture code
**.ends

* expanding   symbol:  double_tail_comp.sym # of pins=10
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/double_tail_comp.sch
.subckt double_tail_comp VDD CLK_bar Vout_n Vout_p Di_p Di_n Vin_n Vin_p CLK VSS
+ Vout_p
X0 VDD.t20 CLK_bar.t0 latch.inv1.VDD VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X1 Vout_p.t5 Vout_n.t8 latch.inv1.VDD VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X2 Di_n.t13 Vin_p.t0 a_88_n1613.t12 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X3 latch.inv1.VDD CLK_bar.t1 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X4 a_88_n1613.t15 Vin_p.t1 Di_n.t12 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X5 VDD.t16 CLK_bar.t2 latch.inv1.VDD VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X6 Vout_p.t1 Di_n.t14 VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X7 a_88_n1613.t23 CLK.t0 VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X8 a_88_n1613.t19 Vin_p.t2 Di_n.t11 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X9 a_88_n1613.t4 Vin_n.t0 Di_p.t13 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X10 VSS.t25 CLK.t1 a_88_n1613.t21 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X11 Di_p.t12 Vin_n.t1 a_88_n1613.t1 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X12 Di_p.t1 CLK.t2 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X13 a_88_n1613.t5 CLK.t3 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X14 VDD.t25 CLK.t4 Di_p.t0 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X15 a_88_n1613.t25 CLK.t5 VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X16 VSS.t51 CLK.t6 a_88_n1613.t32 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X17 a_88_n1613.t18 Vin_p.t3 Di_n.t10 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X18 latch.inv1.VDD Vout_p.t8 Vout_n.t5 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X19 Di_n.t1 CLK.t7 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X20 Vout_n.t1 Vout_p.t9 VSS.t43 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X21 VSS.t30 Di_n.t15 Vout_p.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X22 Di_p.t11 Vin_n.t2 a_88_n1613.t24 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X23 VDD.t2 CLK.t8 Di_n.t0 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X24 a_88_n1613.t29 Vin_n.t3 Di_p.t10 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.81 as=0.237 ps=1.4 w=0.84 l=0.15
X25 latch.inv1.VDD CLK_bar.t3 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X26 VSS.t45 CLK.t9 a_88_n1613.t30 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X27 Di_n.t9 Vin_p.t4 a_88_n1613.t11 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X28 Di_n.t8 Vin_p.t5 a_88_n1613.t8 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X29 Vout_n.t3 Di_p.t14 VSS.t40 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X30 a_88_n1613.t17 Vin_p.t6 Di_n.t7 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X31 a_88_n1613.t10 Vin_p.t7 Di_n.t6 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X32 a_88_n1613.t3 Vin_n.t4 Di_p.t9 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X33 a_88_n1613.t28 Vin_n.t5 Di_p.t8 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X34 Di_n.t5 Vin_p.t8 a_88_n1613.t14 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X35 Di_p.t7 Vin_n.t6 a_88_n1613.t20 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X36 latch.inv1.VDD CLK_bar.t4 VDD.t12 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X37 latch.inv1.VDD Vout_n.t9 Vout_p.t4 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X38 VSS.t42 Vout_p.t10 Vout_n.t7 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X39 Di_p.t6 Vin_n.t7 a_88_n1613.t27 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X40 VDD.t11 CLK_bar.t5 latch.inv1.VDD VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X41 Vout_n.t0 Vout_p.t11 latch.inv1.VDD VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X42 latch.inv1.VDD Vout_p.t12 Vout_n.t4 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X43 a_88_n1613.t33 CLK.t10 VSS.t53 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X44 a_88_n1613.t9 Vin_p.t9 Di_n.t4 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X45 VSS.t47 Di_p.t15 Vout_n.t6 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X46 VSS.t3 CLK.t11 a_88_n1613.t2 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X47 latch.inv1.VDD Vout_n.t10 Vout_p.t3 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X48 Vout_p.t6 Vout_n.t11 VSS.t56 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X49 a_88_n1613.t7 CLK.t12 VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.119 pd=0.985 as=0.121 ps=0.995 w=0.42 l=0.15
X50 Vout_n.t2 Vout_p.t13 latch.inv1.VDD VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X51 VSS.t49 CLK.t13 a_88_n1613.t31 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.121 pd=0.995 as=0.119 ps=0.985 w=0.42 l=0.15
X52 Di_p.t5 Vin_n.t8 a_88_n1613.t22 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.475 ps=2.81 w=0.84 l=0.15
X53 Di_n.t3 Vin_p.t10 a_88_n1613.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X54 a_88_n1613.t6 Vin_n.t9 Di_p.t4 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X55 Vout_p.t2 Vout_n.t12 latch.inv1.VDD VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.119 pd=0.985 as=0.237 ps=1.97 w=0.42 l=0.15
X56 Di_n.t2 Vin_p.t11 a_88_n1613.t16 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
X57 a_88_n1613.t26 Vin_n.t10 Di_p.t3 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.242 pd=1.41 as=0.237 ps=1.4 w=0.84 l=0.15
X58 VSS.t54 Vout_n.t13 Vout_p.t7 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.97 as=0.119 ps=0.985 w=0.42 l=0.15
X59 Di_p.t2 Vin_n.t11 a_88_n1613.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.237 pd=1.4 as=0.242 ps=1.41 w=0.84 l=0.15
R0 CLK_bar.n1 CLK_bar.t3 231.618
R1 CLK_bar.n2 CLK_bar.t1 231.618
R2 CLK_bar.n0 CLK_bar.t4 231.618
R3 CLK_bar.n1 CLK_bar.t0 231.618
R4 CLK_bar.n2 CLK_bar.t5 231.618
R5 CLK_bar.n0 CLK_bar.t2 231.618
R6 CLK_bar CLK_bar.n2 73.9026
R7 CLK_bar CLK_bar.n0 73.9026
R8 CLK_bar CLK_bar.n1 73.311
R9 VDD.n18 VDD.t2 735.818
R10 VDD.n53 VDD.t25 735.818
R11 VDD.n20 VDD.t4 733.472
R12 VDD.n47 VDD.t7 733.472
R13 VDD.n74 VDD.t16 370.702
R14 VDD.n84 VDD.t18 369.529
R15 VDD.n82 VDD.n33 302.69
R16 VDD.n77 VDD.n76 302.69
R17 VDD.n9 VDD.t1 204.514
R18 VDD.n7 VDD.t6 203.571
R19 VDD.n97 VDD.n96 140.934
R20 VDD.n63 VDD.n62 140.934
R21 VDD.n8 VDD.n7 135.714
R22 VDD.n9 VDD.n8 135.714
R23 VDD.t6 VDD.t24 134.773
R24 VDD.t1 VDD.t3 134.773
R25 VDD.n64 VDD.n63 119.71
R26 VDD.n96 VDD.n27 119.71
R27 VDD.n94 VDD.n93 92.5005
R28 VDD.n94 VDD.n27 92.5005
R29 VDD.n95 VDD.n26 92.5005
R30 VDD.n66 VDD.n65 92.5005
R31 VDD.n65 VDD.n64 92.5005
R32 VDD.n44 VDD.n43 92.5005
R33 VDD.n11 VDD.n10 92.5005
R34 VDD.n10 VDD.n9 92.5005
R35 VDD.n3 VDD.n2 92.5005
R36 VDD.n8 VDD.n3 92.5005
R37 VDD.n6 VDD.n5 92.5005
R38 VDD.n7 VDD.n6 92.5005
R39 VDD.n95 VDD.n94 86.4005
R40 VDD.n65 VDD.n44 86.4005
R41 VDD.n6 VDD.n3 86.4005
R42 VDD.n10 VDD.n3 86.4005
R43 VDD.t5 VDD.t15 68.3289
R44 VDD.t9 VDD.t19 68.3289
R45 VDD.n33 VDD.t11 68.0124
R46 VDD.n76 VDD.t20 68.0124
R47 VDD.t13 VDD.t21 67.8576
R48 VDD.t17 VDD.t0 67.8576
R49 VDD.t22 VDD.t5 67.3864
R50 VDD.t15 VDD.t9 67.3864
R51 VDD.t19 VDD.t13 67.3864
R52 VDD.t0 VDD.t8 67.3864
R53 VDD.t10 VDD.t23 66.9152
R54 VDD.n33 VDD.t14 66.8398
R55 VDD.n76 VDD.t12 66.8398
R56 VDD.n64 VDD.t22 34.4003
R57 VDD.t8 VDD.n27 34.4003
R58 VDD.n96 VDD.n95 19.6319
R59 VDD.n63 VDD.n44 19.6319
R60 VDD.n93 VDD.n26 9.2165
R61 VDD.n97 VDD.n26 9.2165
R62 VDD.n62 VDD.n43 9.2165
R63 VDD.n66 VDD.n43 9.2165
R64 VDD.n5 VDD.n2 9.2165
R65 VDD.n11 VDD.n2 9.2165
R66 VDD.n61 VDD.n60 5.12967
R67 VDD.n99 VDD.n98 5.12967
R68 VDD.n92 VDD.n91 5.12967
R69 VDD.n68 VDD.n67 5.12967
R70 VDD.n4 VDD.n0 5.12967
R71 VDD.n13 VDD.n12 5.12967
R72 VDD.n93 VDD.n92 4.6505
R73 VDD.n26 VDD.n25 4.6505
R74 VDD.n98 VDD.n97 4.6505
R75 VDD.n43 VDD.n42 4.6505
R76 VDD.n67 VDD.n66 4.6505
R77 VDD.n62 VDD.n61 4.6505
R78 VDD.n2 VDD.n1 4.6505
R79 VDD.n12 VDD.n11 4.6505
R80 VDD.n5 VDD.n4 4.6505
R81 VDD.n59 VDD.n56 3.43958
R82 VDD.n101 VDD.n100 3.43958
R83 VDD.n55 VDD.n54 3.43958
R84 VDD.n102 VDD.n21 3.43958
R85 VDD.n30 VDD.n24 3.4105
R86 VDD.n41 VDD.n40 3.4105
R87 VDD.n69 VDD.n68 3.4105
R88 VDD.n38 VDD.n37 3.4105
R89 VDD.n74 VDD.n73 3.4105
R90 VDD.n75 VDD.n36 3.4105
R91 VDD.n78 VDD.n77 3.4105
R92 VDD.n34 VDD 3.4105
R93 VDD.n82 VDD.n81 3.4105
R94 VDD.n83 VDD.n32 3.4105
R95 VDD.n85 VDD.n84 3.4105
R96 VDD.n29 VDD.n28 3.4105
R97 VDD.n91 VDD.n90 3.4105
R98 VDD.n52 VDD.n51 3.4105
R99 VDD.n48 VDD.n47 3.4105
R100 VDD.n14 VDD.n0 3.4105
R101 VDD VDD.n110 3.4105
R102 VDD.n15 VDD.n13 3.4105
R103 VDD.n106 VDD.n18 3.4105
R104 VDD.n105 VDD.n19 3.4105
R105 VDD.n46 VDD.n45 3.4105
R106 VDD.n51 VDD.n50 3.4105
R107 VDD.n49 VDD.n48 3.4105
R108 VDD.n16 VDD.n14 3.4105
R109 VDD.n110 VDD.n109 3.4105
R110 VDD.n108 VDD.n15 3.4105
R111 VDD.n107 VDD.n106 3.4105
R112 VDD.n105 VDD.n17 3.4105
R113 VDD.n104 VDD.n103 3.4105
R114 VDD.n88 VDD.n30 3.4105
R115 VDD.n23 VDD.n22 3.4105
R116 VDD.n58 VDD.n57 3.4105
R117 VDD.n40 VDD.n39 3.4105
R118 VDD.n70 VDD.n69 3.4105
R119 VDD.n71 VDD.n38 3.4105
R120 VDD.n73 VDD.n72 3.4105
R121 VDD.n36 VDD.n35 3.4105
R122 VDD.n79 VDD.n78 3.4105
R123 VDD VDD.n34 3.4105
R124 VDD.n81 VDD.n80 3.4105
R125 VDD.n32 VDD.n31 3.4105
R126 VDD.n86 VDD.n85 3.4105
R127 VDD.n87 VDD.n29 3.4105
R128 VDD.n90 VDD.n89 3.4105
R129 VDD.n102 VDD.n101 1.93491
R130 VDD.n56 VDD.n55 1.93491
R131 VDD.n60 VDD.n59 1.72871
R132 VDD.n100 VDD.n99 1.72871
R133 VDD.n54 VDD.n53 1.72871
R134 VDD.n21 VDD.n20 1.72871
R135 VDD.t21 VDD.t10 0.47173
R136 VDD.t23 VDD.t17 0.47173
R137 VDD.n60 VDD.n41 0.1505
R138 VDD.n68 VDD.n41 0.1505
R139 VDD.n68 VDD.n37 0.1505
R140 VDD.n74 VDD.n37 0.1505
R141 VDD.n75 VDD.n74 0.1505
R142 VDD.n77 VDD.n75 0.1505
R143 VDD.n77 VDD 0.1505
R144 VDD.n82 VDD 0.1505
R145 VDD.n83 VDD.n82 0.1505
R146 VDD.n84 VDD.n83 0.1505
R147 VDD.n84 VDD.n28 0.1505
R148 VDD.n91 VDD.n28 0.1505
R149 VDD.n91 VDD.n24 0.1505
R150 VDD.n99 VDD.n24 0.1505
R151 VDD.n53 VDD.n52 0.1505
R152 VDD.n52 VDD.n47 0.1505
R153 VDD.n47 VDD.n0 0.1505
R154 VDD VDD.n0 0.1505
R155 VDD VDD.n13 0.1505
R156 VDD.n18 VDD.n13 0.1505
R157 VDD.n19 VDD.n18 0.1505
R158 VDD.n20 VDD.n19 0.1505
R159 VDD.n92 VDD.n25 0.0905
R160 VDD.n98 VDD.n25 0.0905
R161 VDD.n61 VDD.n42 0.0905
R162 VDD.n67 VDD.n42 0.0905
R163 VDD.n4 VDD.n1 0.0905
R164 VDD.n12 VDD.n1 0.0905
R165 VDD.n58 VDD.n40 0.0569
R166 VDD.n69 VDD.n40 0.0569
R167 VDD.n69 VDD.n38 0.0569
R168 VDD.n73 VDD.n38 0.0569
R169 VDD.n73 VDD.n36 0.0569
R170 VDD.n78 VDD.n36 0.0569
R171 VDD.n78 VDD.n34 0.0569
R172 VDD.n81 VDD.n34 0.0569
R173 VDD.n81 VDD.n32 0.0569
R174 VDD.n85 VDD.n32 0.0569
R175 VDD.n85 VDD.n29 0.0569
R176 VDD.n90 VDD.n29 0.0569
R177 VDD.n90 VDD.n30 0.0569
R178 VDD.n30 VDD.n23 0.0569
R179 VDD.n51 VDD.n46 0.0569
R180 VDD.n51 VDD.n48 0.0569
R181 VDD.n48 VDD.n14 0.0569
R182 VDD.n110 VDD.n14 0.0569
R183 VDD.n110 VDD.n15 0.0569
R184 VDD.n106 VDD.n15 0.0569
R185 VDD.n106 VDD.n105 0.0569
R186 VDD.n105 VDD.n104 0.0569
R187 VDD.n55 VDD.n45 0.03434
R188 VDD.n50 VDD.n45 0.03434
R189 VDD.n50 VDD.n49 0.03434
R190 VDD.n49 VDD.n16 0.03434
R191 VDD.n109 VDD.n16 0.03434
R192 VDD.n109 VDD.n108 0.03434
R193 VDD.n108 VDD.n107 0.03434
R194 VDD.n107 VDD.n17 0.03434
R195 VDD.n103 VDD.n17 0.03434
R196 VDD.n103 VDD.n102 0.03434
R197 VDD.n57 VDD.n56 0.03434
R198 VDD.n57 VDD.n39 0.03434
R199 VDD.n70 VDD.n39 0.03434
R200 VDD.n71 VDD.n70 0.03434
R201 VDD.n72 VDD.n71 0.03434
R202 VDD.n72 VDD.n35 0.03434
R203 VDD.n79 VDD.n35 0.03434
R204 VDD VDD.n79 0.03434
R205 VDD.n80 VDD 0.03434
R206 VDD.n80 VDD.n31 0.03434
R207 VDD.n86 VDD.n31 0.03434
R208 VDD.n87 VDD.n86 0.03434
R209 VDD.n89 VDD.n87 0.03434
R210 VDD.n89 VDD.n88 0.03434
R211 VDD.n88 VDD.n22 0.03434
R212 VDD.n101 VDD.n22 0.03434
R213 VDD.n100 VDD.n23 0.0283716
R214 VDD.n59 VDD.n58 0.0283716
R215 VDD.n54 VDD.n46 0.0283716
R216 VDD.n104 VDD.n21 0.0283716
R217 Vout_n.n2 Vout_n.n1 599.173
R218 Vout_n.n2 Vout_n.n0 599.173
R219 Vout_n.n11 Vout_n.n9 200.374
R220 Vout_n.n11 Vout_n.n10 198.894
R221 Vout_n.n3 Vout_n.t9 164.137
R222 Vout_n.n3 Vout_n.t8 164.137
R223 Vout_n.n4 Vout_n.t10 164.137
R224 Vout_n.n4 Vout_n.t12 164.137
R225 Vout_n.n6 Vout_n.t11 164.137
R226 Vout_n.n6 Vout_n.t13 164.137
R227 Vout_n.n1 Vout_n.t2 133.679
R228 Vout_n.n0 Vout_n.t0 133.679
R229 Vout_n.n1 Vout_n.t5 131.333
R230 Vout_n.n0 Vout_n.t4 131.333
R231 Vout_n.n10 Vout_n.t1 81.4291
R232 Vout_n.n9 Vout_n.t3 81.4291
R233 Vout_n.n10 Vout_n.t7 80.0005
R234 Vout_n.n9 Vout_n.t6 80.0005
R235 Vout_n Vout_n.n6 77.2722
R236 Vout_n.n5 Vout_n.n4 73.9428
R237 Vout_n.n5 Vout_n.n3 73.3637
R238 Vout_n Vout_n.n7 4.14383
R239 Vout_n.n8 Vout_n 4.14383
R240 Vout_n Vout_n.n11 3.85543
R241 Vout_n.n8 Vout_n.n2 3.73637
R242 Vout_n.n7 Vout_n.n5 3.51077
R243 Vout_n.n7 Vout_n 0.107033
R244 Vout_n Vout_n.n8 0.107033
R245 Vout_p.n6 Vout_p.n5 599.173
R246 Vout_p.n6 Vout_p.n4 599.173
R247 Vout_p.n9 Vout_p.n8 200.374
R248 Vout_p.n9 Vout_p.n7 198.894
R249 Vout_p.n1 Vout_p.t8 164.137
R250 Vout_p.n1 Vout_p.t13 164.137
R251 Vout_p.n0 Vout_p.t12 164.137
R252 Vout_p.n0 Vout_p.t11 164.137
R253 Vout_p.n3 Vout_p.t9 164.137
R254 Vout_p.n3 Vout_p.t10 164.137
R255 Vout_p.n5 Vout_p.t3 133.679
R256 Vout_p.n4 Vout_p.t4 133.679
R257 Vout_p.n5 Vout_p.t2 131.333
R258 Vout_p.n4 Vout_p.t5 131.333
R259 Vout_p.n7 Vout_p.t7 81.4291
R260 Vout_p.n8 Vout_p.t1 81.4291
R261 Vout_p.n7 Vout_p.t6 80.0005
R262 Vout_p.n8 Vout_p.t0 80.0005
R263 Vout_p.n11 Vout_p.n3 77.1531
R264 Vout_p.n2 Vout_p.n0 73.9428
R265 Vout_p.n2 Vout_p.n1 73.3637
R266 Vout_p Vout_p.n10 4.14383
R267 Vout_p.n11 Vout_p 4.14383
R268 Vout_p Vout_p.n6 3.85543
R269 Vout_p.n10 Vout_p.n9 3.73637
R270 Vout_p Vout_p.n2 3.62983
R271 Vout_p.n10 Vout_p 0.107033
R272 Vout_p Vout_p.n11 0.107033
R273 Vin_p.n8 Vin_p.t8 231.618
R274 Vin_p.n6 Vin_p.t11 231.618
R275 Vin_p.n5 Vin_p.t4 231.618
R276 Vin_p.n3 Vin_p.t10 231.618
R277 Vin_p.n1 Vin_p.t5 231.618
R278 Vin_p.n0 Vin_p.t0 231.618
R279 Vin_p.n8 Vin_p.t9 231.618
R280 Vin_p.n6 Vin_p.t2 231.618
R281 Vin_p.n5 Vin_p.t6 231.618
R282 Vin_p.n3 Vin_p.t3 231.618
R283 Vin_p.n1 Vin_p.t7 231.618
R284 Vin_p.n0 Vin_p.t1 231.618
R285 Vin_p.n7 Vin_p.n5 73.9026
R286 Vin_p.n2 Vin_p.n0 73.9026
R287 Vin_p.n9 Vin_p.n8 73.311
R288 Vin_p.n7 Vin_p.n6 73.311
R289 Vin_p.n4 Vin_p.n3 73.311
R290 Vin_p.n2 Vin_p.n1 73.311
R291 Vin_p.n9 Vin_p.n7 0.592167
R292 Vin_p.n4 Vin_p.n2 0.592167
R293 Vin_p Vin_p.n9 0.296333
R294 Vin_p Vin_p.n4 0.296333
R295 a_88_n1613.n3 a_88_n1613.n16 198.894
R296 a_88_n1613.n3 a_88_n1613.n15 198.894
R297 a_88_n1613.n2 a_88_n1613.n14 198.894
R298 a_88_n1613.n2 a_88_n1613.n13 198.894
R299 a_88_n1613.n2 a_88_n1613.n12 198.894
R300 a_88_n1613.n1 a_88_n1613.t15 144.418
R301 a_88_n1613.n0 a_88_n1613.t29 144.418
R302 a_88_n1613.n1 a_88_n1613.t11 143.703
R303 a_88_n1613.n0 a_88_n1613.t22 143.703
R304 a_88_n1613.t28 a_88_n1613.n0 102.689
R305 a_88_n1613.n1 a_88_n1613.n9 102.689
R306 a_88_n1613.n1 a_88_n1613.n10 102.689
R307 a_88_n1613.n1 a_88_n1613.n11 102.689
R308 a_88_n1613.n1 a_88_n1613.n8 102.689
R309 a_88_n1613.n1 a_88_n1613.n7 102.689
R310 a_88_n1613.n0 a_88_n1613.n5 102.689
R311 a_88_n1613.n0 a_88_n1613.n6 102.689
R312 a_88_n1613.n0 a_88_n1613.n17 102.689
R313 a_88_n1613.n0 a_88_n1613.n4 102.689
R314 a_88_n1613.n16 a_88_n1613.t23 81.4291
R315 a_88_n1613.n15 a_88_n1613.t25 81.4291
R316 a_88_n1613.n14 a_88_n1613.t5 81.4291
R317 a_88_n1613.n13 a_88_n1613.t7 81.4291
R318 a_88_n1613.n12 a_88_n1613.t33 81.4291
R319 a_88_n1613.n16 a_88_n1613.t21 80.0005
R320 a_88_n1613.n15 a_88_n1613.t31 80.0005
R321 a_88_n1613.n14 a_88_n1613.t2 80.0005
R322 a_88_n1613.n13 a_88_n1613.t32 80.0005
R323 a_88_n1613.n12 a_88_n1613.t30 80.0005
R324 a_88_n1613.n9 a_88_n1613.t17 41.4291
R325 a_88_n1613.n10 a_88_n1613.t19 41.4291
R326 a_88_n1613.n11 a_88_n1613.t9 41.4291
R327 a_88_n1613.n8 a_88_n1613.t18 41.4291
R328 a_88_n1613.n7 a_88_n1613.t10 41.4291
R329 a_88_n1613.n5 a_88_n1613.t6 41.4291
R330 a_88_n1613.n6 a_88_n1613.t3 41.4291
R331 a_88_n1613.n17 a_88_n1613.t26 41.4291
R332 a_88_n1613.n4 a_88_n1613.t4 41.4291
R333 a_88_n1613.n9 a_88_n1613.t16 40.7148
R334 a_88_n1613.n10 a_88_n1613.t14 40.7148
R335 a_88_n1613.n11 a_88_n1613.t13 40.7148
R336 a_88_n1613.n8 a_88_n1613.t8 40.7148
R337 a_88_n1613.n7 a_88_n1613.t12 40.7148
R338 a_88_n1613.n5 a_88_n1613.t1 40.7148
R339 a_88_n1613.n6 a_88_n1613.t27 40.7148
R340 a_88_n1613.n17 a_88_n1613.t24 40.7148
R341 a_88_n1613.n4 a_88_n1613.t20 40.7148
R342 a_88_n1613.t0 a_88_n1613.t28 40.7148
R343 a_88_n1613.n2 a_88_n1613.n1 12.2838
R344 a_88_n1613.n0 a_88_n1613.n3 12.2838
R345 a_88_n1613.n3 a_88_n1613.n2 2.36717
R346 Di_n Di_n.n1 603.328
R347 Di_n.n0 Di_n.t15 164.137
R348 Di_n.n0 Di_n.t14 164.137
R349 Di_n.n1 Di_n.t1 133.679
R350 Di_n.n1 Di_n.t0 131.333
R351 Di_n.n10 Di_n.n8 102.382
R352 Di_n.n3 Di_n.n2 101.79
R353 Di_n.n5 Di_n.n4 101.79
R354 Di_n.n7 Di_n.n6 101.79
R355 Di_n.n12 Di_n.n11 101.79
R356 Di_n.n10 Di_n.n9 101.79
R357 Di_n Di_n.n0 73.3637
R358 Di_n.n2 Di_n.t13 40.7148
R359 Di_n.n4 Di_n.t8 40.7148
R360 Di_n.n6 Di_n.t3 40.7148
R361 Di_n.n11 Di_n.t5 40.7148
R362 Di_n.n9 Di_n.t2 40.7148
R363 Di_n.n8 Di_n.t9 40.7148
R364 Di_n.n2 Di_n.t12 40.0005
R365 Di_n.n4 Di_n.t6 40.0005
R366 Di_n.n6 Di_n.t10 40.0005
R367 Di_n.n11 Di_n.t4 40.0005
R368 Di_n.n9 Di_n.t11 40.0005
R369 Di_n.n8 Di_n.t7 40.0005
R370 Di_n Di_n.n13 8.49997
R371 Di_n.n3 Di_n 4.4346
R372 Di_n.n12 Di_n.n10 0.592167
R373 Di_n.n7 Di_n.n5 0.592167
R374 Di_n.n5 Di_n.n3 0.592167
R375 Di_n.n13 Di_n.n12 0.279667
R376 Di_n.n13 Di_n.n7 0.279667
R377 VSS.n53 VSS.n52 63308.6
R378 VSS.n51 VSS.n19 37145.5
R379 VSS.n60 VSS.n18 585
R380 VSS.n66 VSS.n18 585
R381 VSS.n17 VSS.n16 585
R382 VSS.n67 VSS.n17 585
R383 VSS.n70 VSS.n69 585
R384 VSS.n69 VSS.n68 585
R385 VSS.n49 VSS.n48 585
R386 VSS.n50 VSS.n49 585
R387 VSS.n25 VSS.n24 585
R388 VSS.n24 VSS.n22 585
R389 VSS.n44 VSS.n43 585
R390 VSS.n43 VSS.n42 585
R391 VSS.n65 VSS.n64 585
R392 VSS.n66 VSS.n65 585
R393 VSS.n21 VSS.n20 585
R394 VSS.n54 VSS.n20 585
R395 VSS.n57 VSS.n56 585
R396 VSS.n56 VSS.n55 585
R397 VSS.n37 VSS.n36 585
R398 VSS.n36 VSS.n35 585
R399 VSS.n33 VSS.n32 585
R400 VSS.n34 VSS.n33 585
R401 VSS.n31 VSS.n23 585
R402 VSS.n50 VSS.n23 585
R403 VSS.n74 VSS.t30 282.651
R404 VSS.n76 VSS.t56 282.651
R405 VSS.n0 VSS.t42 282.651
R406 VSS.n27 VSS.t25 282.651
R407 VSS.n75 VSS.t53 281.223
R408 VSS.n12 VSS.t54 281.223
R409 VSS.n2 VSS.t43 281.223
R410 VSS.n28 VSS.t40 281.223
R411 VSS.n39 VSS.t47 278.151
R412 VSS.n72 VSS.t32 276.723
R413 VSS.t37 VSS.t4 210.98
R414 VSS.t34 VSS.t2 210.98
R415 VSS.t6 VSS.t50 210.98
R416 VSS.t17 VSS.t19 210.98
R417 VSS.t46 VSS.t39 208.07
R418 VSS.t36 VSS.t37 208.07
R419 VSS.t4 VSS.t1 208.07
R420 VSS.t24 VSS.t27 208.07
R421 VSS.t8 VSS.t26 208.07
R422 VSS.t48 VSS.t34 208.07
R423 VSS.t2 VSS.t6 208.07
R424 VSS.t50 VSS.t9 208.07
R425 VSS.t44 VSS.t52 208.07
R426 VSS.t15 VSS.t17 208.07
R427 VSS.t19 VSS.t12 208.07
R428 VSS.t29 VSS.t31 208.07
R429 VSS.t21 VSS.t55 206.614
R430 VSS VSS.n13 199.794
R431 VSS.n9 VSS.n8 199.794
R432 VSS.n7 VSS.n6 199.794
R433 VSS VSS.n1 199.794
R434 VSS.n65 VSS.n20 164.93
R435 VSS.n56 VSS.n20 164.93
R436 VSS.n43 VSS.n24 164.93
R437 VSS.n49 VSS.n24 164.93
R438 VSS.n69 VSS.n17 164.93
R439 VSS.n18 VSS.n17 164.93
R440 VSS.n33 VSS.n23 164.93
R441 VSS.n36 VSS.n33 164.93
R442 VSS.t38 VSS.n34 106.218
R443 VSS.n67 VSS.t20 106.218
R444 VSS.t16 VSS.n54 106.218
R445 VSS.n42 VSS.t23 104.763
R446 VSS.t23 VSS.n22 104.763
R447 VSS.n50 VSS.t0 104.763
R448 VSS.n34 VSS.t0 104.763
R449 VSS.n35 VSS.t33 104.763
R450 VSS.n68 VSS.t14 104.763
R451 VSS.t14 VSS.n67 104.763
R452 VSS.n55 VSS.t18 104.763
R453 VSS.n42 VSS.t41 103.308
R454 VSS.n35 VSS.t38 103.308
R455 VSS.n68 VSS.t13 103.308
R456 VSS.t20 VSS.n66 103.308
R457 VSS.n55 VSS.t16 103.308
R458 VSS.n13 VSS.t45 82.8576
R459 VSS.n8 VSS.t51 82.8576
R460 VSS.n6 VSS.t3 82.8576
R461 VSS.n1 VSS.t49 82.8576
R462 VSS.n13 VSS.t10 81.4291
R463 VSS.n8 VSS.t7 81.4291
R464 VSS.n6 VSS.t35 81.4291
R465 VSS.n1 VSS.t28 81.4291
R466 VSS.n52 VSS.n22 64.0217
R467 VSS.t11 VSS.n19 64.0217
R468 VSS.n54 VSS.n53 64.0217
R469 VSS.t5 VSS.n51 62.5666
R470 VSS.n52 VSS.t5 42.1963
R471 VSS.n51 VSS.n50 40.7412
R472 VSS.n66 VSS.n19 40.7412
R473 VSS.n53 VSS.t11 40.7412
R474 VSS.n44 VSS.n25 10.7168
R475 VSS.n48 VSS.n25 10.7168
R476 VSS.n64 VSS.n21 10.7168
R477 VSS.n57 VSS.n21 10.7168
R478 VSS.n70 VSS.n16 10.7168
R479 VSS.n60 VSS.n16 10.7168
R480 VSS.n32 VSS.n31 10.7168
R481 VSS.n37 VSS.n32 10.7168
R482 VSS.n46 VSS.n25 9.3005
R483 VSS.n48 VSS.n47 9.3005
R484 VSS.n45 VSS.n44 9.3005
R485 VSS.n64 VSS.n63 9.3005
R486 VSS.n59 VSS.n21 9.3005
R487 VSS.n58 VSS.n57 9.3005
R488 VSS.n16 VSS.n15 9.3005
R489 VSS.n61 VSS.n60 9.3005
R490 VSS.n71 VSS.n70 9.3005
R491 VSS.n32 VSS.n29 9.3005
R492 VSS.n38 VSS.n37 9.3005
R493 VSS.n31 VSS.n30 9.3005
R494 VSS.n45 VSS.n41 5.71717
R495 VSS.n58 VSS.n14 5.71717
R496 VSS.n41 VSS.n26 4.5005
R497 VSS.n40 VSS.n39 4.5005
R498 VSS.n62 VSS.n14 4.5005
R499 VSS.n73 VSS.n72 4.5005
R500 VSS.n75 VSS.n11 3.43911
R501 VSS.n27 VSS.n5 3.43911
R502 VSS.n3 VSS.n0 3.4105
R503 VSS VSS.n88 3.4105
R504 VSS.n4 VSS.n2 3.4105
R505 VSS.n84 VSS.n7 3.4105
R506 VSS.n83 VSS 3.4105
R507 VSS.n82 VSS.n9 3.4105
R508 VSS.n12 VSS.n10 3.4105
R509 VSS.n78 VSS 3.4105
R510 VSS.n77 VSS.n76 3.4105
R511 VSS.n88 VSS.n87 3.4105
R512 VSS.n86 VSS.n4 3.4105
R513 VSS.n85 VSS.n84 3.4105
R514 VSS.n83 VSS 3.4105
R515 VSS.n82 VSS.n81 3.4105
R516 VSS.n80 VSS.n10 3.4105
R517 VSS.n79 VSS.n78 3.4105
R518 VSS.n87 VSS.n5 1.73427
R519 VSS.n79 VSS.n11 1.73427
R520 VSS.t33 VSS.t46 1.45553
R521 VSS.t39 VSS.t36 1.45553
R522 VSS.t1 VSS.t24 1.45553
R523 VSS.t27 VSS.t8 1.45553
R524 VSS.t26 VSS.t48 1.45553
R525 VSS.t9 VSS.t21 1.45553
R526 VSS.t55 VSS.t22 1.45553
R527 VSS.t22 VSS.t44 1.45553
R528 VSS.t52 VSS.t15 1.45553
R529 VSS.t12 VSS.t29 1.45553
R530 VSS.t31 VSS.t13 1.45553
R531 VSS.n39 VSS.n38 0.917167
R532 VSS.n47 VSS.n26 0.917167
R533 VSS.n72 VSS.n71 0.917167
R534 VSS.n63 VSS.n62 0.917167
R535 VSS.n62 VSS.n61 0.917167
R536 VSS.n30 VSS.n26 0.917167
R537 VSS.n41 VSS.n40 0.3005
R538 VSS.n40 VSS.n28 0.3005
R539 VSS.n28 VSS.n27 0.3005
R540 VSS.n75 VSS.n74 0.3005
R541 VSS.n74 VSS.n73 0.3005
R542 VSS.n73 VSS.n14 0.3005
R543 VSS.n27 VSS.n0 0.1505
R544 VSS VSS.n0 0.1505
R545 VSS VSS.n2 0.1505
R546 VSS.n7 VSS.n2 0.1505
R547 VSS VSS.n7 0.1505
R548 VSS.n9 VSS 0.1505
R549 VSS.n12 VSS.n9 0.1505
R550 VSS VSS.n12 0.1505
R551 VSS.n76 VSS 0.1505
R552 VSS.n76 VSS.n75 0.1505
R553 VSS.n46 VSS.n45 0.105151
R554 VSS.n47 VSS.n46 0.105151
R555 VSS.n63 VSS.n59 0.105151
R556 VSS.n59 VSS.n58 0.105151
R557 VSS.n71 VSS.n15 0.105151
R558 VSS.n61 VSS.n15 0.105151
R559 VSS.n30 VSS.n29 0.105151
R560 VSS.n38 VSS.n29 0.105151
R561 VSS.n88 VSS.n3 0.0569
R562 VSS.n88 VSS.n4 0.0569
R563 VSS.n84 VSS.n4 0.0569
R564 VSS.n84 VSS.n83 0.0569
R565 VSS.n83 VSS.n82 0.0569
R566 VSS.n82 VSS.n10 0.0569
R567 VSS.n78 VSS.n10 0.0569
R568 VSS.n78 VSS.n77 0.0569
R569 VSS.n87 VSS.n86 0.03434
R570 VSS.n86 VSS.n85 0.03434
R571 VSS.n85 VSS 0.03434
R572 VSS.n81 VSS 0.03434
R573 VSS.n81 VSS.n80 0.03434
R574 VSS.n80 VSS.n79 0.03434
R575 VSS.n5 VSS.n3 0.0288317
R576 VSS.n77 VSS.n11 0.0288317
R577 CLK.n3 CLK.t11 164.137
R578 CLK.n3 CLK.t3 164.137
R579 CLK.n8 CLK.t7 164.137
R580 CLK.n8 CLK.t8 164.137
R581 CLK.n7 CLK.t2 164.137
R582 CLK.n7 CLK.t4 164.137
R583 CLK.n5 CLK.t6 164.137
R584 CLK.n5 CLK.t12 164.137
R585 CLK.n4 CLK.t9 164.137
R586 CLK.n4 CLK.t10 164.137
R587 CLK.n1 CLK.t13 164.137
R588 CLK.n1 CLK.t5 164.137
R589 CLK.n0 CLK.t1 164.137
R590 CLK.n0 CLK.t0 164.137
R591 CLK.n9 CLK.n8 74.2428
R592 CLK.n9 CLK.n7 74.2428
R593 CLK.n6 CLK.n4 73.9553
R594 CLK.n2 CLK.n0 73.9553
R595 CLK CLK.n3 73.3637
R596 CLK.n6 CLK.n5 73.3637
R597 CLK.n2 CLK.n1 73.3637
R598 CLK CLK.n9 8.04877
R599 CLK CLK.n6 0.579667
R600 CLK CLK.n2 0.579667
R601 Vin_n.n8 Vin_n.t7 231.618
R602 Vin_n.n6 Vin_n.t1 231.618
R603 Vin_n.n5 Vin_n.t8 231.618
R604 Vin_n.n3 Vin_n.t2 231.618
R605 Vin_n.n1 Vin_n.t11 231.618
R606 Vin_n.n0 Vin_n.t6 231.618
R607 Vin_n.n8 Vin_n.t10 231.618
R608 Vin_n.n6 Vin_n.t4 231.618
R609 Vin_n.n5 Vin_n.t9 231.618
R610 Vin_n.n3 Vin_n.t5 231.618
R611 Vin_n.n1 Vin_n.t0 231.618
R612 Vin_n.n0 Vin_n.t3 231.618
R613 Vin_n.n7 Vin_n.n5 73.9026
R614 Vin_n.n2 Vin_n.n0 73.9026
R615 Vin_n.n9 Vin_n.n8 73.311
R616 Vin_n.n7 Vin_n.n6 73.311
R617 Vin_n.n4 Vin_n.n3 73.311
R618 Vin_n.n2 Vin_n.n1 73.311
R619 Vin_n.n9 Vin_n.n7 0.592167
R620 Vin_n.n4 Vin_n.n2 0.592167
R621 Vin_n Vin_n.n9 0.296333
R622 Vin_n Vin_n.n4 0.296333
R623 Di_p Di_p.n6 603.328
R624 Di_p.n0 Di_p.t15 164.137
R625 Di_p.n0 Di_p.t14 164.137
R626 Di_p.n6 Di_p.t1 133.679
R627 Di_p.n6 Di_p.t0 131.333
R628 Di_p.n3 Di_p.n1 102.382
R629 Di_p.n8 Di_p.n7 101.79
R630 Di_p.n10 Di_p.n9 101.79
R631 Di_p.n12 Di_p.n11 101.79
R632 Di_p.n5 Di_p.n4 101.79
R633 Di_p.n3 Di_p.n2 101.79
R634 Di_p Di_p.n0 73.3637
R635 Di_p.n7 Di_p.t5 40.7148
R636 Di_p.n9 Di_p.t12 40.7148
R637 Di_p.n11 Di_p.t6 40.7148
R638 Di_p.n4 Di_p.t11 40.7148
R639 Di_p.n2 Di_p.t2 40.7148
R640 Di_p.n1 Di_p.t7 40.7148
R641 Di_p.n7 Di_p.t4 40.0005
R642 Di_p.n9 Di_p.t9 40.0005
R643 Di_p.n11 Di_p.t3 40.0005
R644 Di_p.n4 Di_p.t8 40.0005
R645 Di_p.n2 Di_p.t13 40.0005
R646 Di_p.n1 Di_p.t10 40.0005
R647 Di_p Di_p.n13 8.49997
R648 Di_p.n8 Di_p 4.4346
R649 Di_p.n5 Di_p.n3 0.592167
R650 Di_p.n12 Di_p.n10 0.592167
R651 Di_p.n10 Di_p.n8 0.592167
R652 Di_p.n13 Di_p.n5 0.279667
R653 Di_p.n13 Di_p.n12 0.279667
C0 latch.inv1.VDD VDD 2.82f
.ends



* expanding   symbol:  RS_latch.sym # of pins=5
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/RS_latch.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/RS_latch.sch
.subckt RS_latch VDD R Q S Q_bar
*.iopin VDD
*.opin Q
*.opin Q_bar
*.ipin R
*.ipin S
x1 VDD R Q_bar Q nor
x2 VDD Q S Q_bar nor
.ends


* expanding   symbol:  nor.sym # of pins=4
** sym_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/nor.sym
** sch_path: /fs1/eecg/tcc/lizongh2/sky130_comparator/xschem/nor.sch
.subckt nor VDD A B out
*.iopin VDD
*.ipin A
*.ipin B
*.opin out
XM1 out B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 out B net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
**** begin user architecture code

.model filesrc filesource (file="staircase_voltage.txt" amploffset=[Vcm] amplscale=[1] timeoffset=0
+ timescale=1 timerelative=false amplstep=false)

**** end user architecture code
.end

magic
tech sky130A
magscale 1 2
timestamp 1706046249
<< nwell >>
rect -36 -42 292 210
<< pmos >>
rect 113 0 143 168
<< pdiff >>
rect 0 146 113 168
rect 0 106 36 146
rect 76 106 113 146
rect 0 62 113 106
rect 0 22 36 62
rect 76 22 113 62
rect 0 0 113 22
rect 143 146 256 168
rect 143 106 180 146
rect 220 106 256 146
rect 143 62 256 106
rect 143 22 180 62
rect 220 22 256 62
rect 143 0 256 22
<< pdiffc >>
rect 36 106 76 146
rect 36 22 76 62
rect 180 106 220 146
rect 180 22 220 62
<< poly >>
rect 88 264 168 284
rect 88 224 108 264
rect 148 224 168 264
rect 88 204 168 224
rect 113 168 143 204
rect 113 -36 143 0
<< polycont >>
rect 108 224 148 264
<< locali >>
rect 88 264 168 284
rect 88 224 108 264
rect 148 224 168 264
rect 88 204 168 224
rect 26 146 86 162
rect 26 106 36 146
rect 76 106 86 146
rect 26 62 86 106
rect 26 22 36 62
rect 76 22 86 62
rect 26 6 86 22
rect 170 146 230 162
rect 170 106 180 146
rect 220 106 230 146
rect 170 62 230 106
rect 170 22 180 62
rect 220 22 230 62
rect 170 6 230 22
<< viali >>
rect 108 224 148 264
rect 36 106 76 146
rect 36 22 76 62
rect 180 106 220 146
rect 180 22 220 62
<< metal1 >>
rect 88 264 168 284
rect 88 224 108 264
rect 148 224 168 264
rect 88 204 168 224
rect 26 146 86 162
rect 26 106 36 146
rect 76 106 86 146
rect 26 62 86 106
rect 26 22 36 62
rect 76 22 86 62
rect 26 -42 86 22
rect 170 146 230 162
rect 170 106 180 146
rect 220 106 230 146
rect 170 62 230 106
rect 170 22 180 62
rect 220 22 230 62
rect 170 -42 230 22
<< end >>

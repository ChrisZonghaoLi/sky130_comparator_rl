.param Vcm=0.9008961886167527
.param VDD=1.8
.param Vin=0.05
.param Vin_min=0.0001
.param CL=2e-14
.param Tclk=1e-09
.param Tclk_pk=4.5e-10
.param Tdelay=2e-10
.param Tdelay_bar=7.000000000000001e-10
.param Tr=5.000000000000001e-11
.param Tf=5.000000000000001e-11
  
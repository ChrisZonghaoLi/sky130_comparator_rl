* NGSPICE file created from nfet_01v8_0p84_nf1.ext - technology: sky130A

.subckt nfet_01v8_0p84_nf1
X0 a_143_0# a_88_204# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.81 as=0.475 ps=2.81 w=0.84 l=0.15
.ends

